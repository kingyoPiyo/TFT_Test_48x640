/***********************************************************************************
* Title    : 🍣 ROM
* Date     : 2021/01/11
* Design   : kingyo
* Note     : 🍣 data from : https://github.com/htlabnet/inside_magimajopures
***********************************************************************************/
module sushi_rom (
    input   wire            i_clk,
    input   wire    [11:0]  i_addr,
    output  reg     [15:0]  o_data
    )/* synthesis syn_romstyle = "block_rom" */;

    always @(posedge i_clk) begin
        case (i_addr[11:0])
            12'd0 : o_data <= 16'h0000;
            12'd1 : o_data <= 16'h0000;
            12'd2 : o_data <= 16'h0000;
            12'd3 : o_data <= 16'h0000;
            12'd4 : o_data <= 16'h0000;
            12'd5 : o_data <= 16'h0000;
            12'd6 : o_data <= 16'h0000;
            12'd7 : o_data <= 16'h0000;
            12'd8 : o_data <= 16'h0000;
            12'd9 : o_data <= 16'h0000;
            12'd10 : o_data <= 16'h0000;
            12'd11 : o_data <= 16'h0000;
            12'd12 : o_data <= 16'h0000;
            12'd13 : o_data <= 16'h0000;
            12'd14 : o_data <= 16'h0000;
            12'd15 : o_data <= 16'h0000;
            12'd16 : o_data <= 16'h0000;
            12'd17 : o_data <= 16'h0000;
            12'd18 : o_data <= 16'h0000;
            12'd19 : o_data <= 16'h0000;
            12'd20 : o_data <= 16'h0000;
            12'd21 : o_data <= 16'h0000;
            12'd22 : o_data <= 16'h0000;
            12'd23 : o_data <= 16'h0000;
            12'd24 : o_data <= 16'h0000;
            12'd25 : o_data <= 16'h0000;
            12'd26 : o_data <= 16'h0000;
            12'd27 : o_data <= 16'h0000;
            12'd28 : o_data <= 16'h0000;
            12'd29 : o_data <= 16'h0000;
            12'd30 : o_data <= 16'h0000;
            12'd31 : o_data <= 16'h0000;
            12'd32 : o_data <= 16'h0000;
            12'd33 : o_data <= 16'h0000;
            12'd34 : o_data <= 16'h0000;
            12'd35 : o_data <= 16'h0000;
            12'd36 : o_data <= 16'h0000;
            12'd37 : o_data <= 16'h0000;
            12'd38 : o_data <= 16'h0000;
            12'd39 : o_data <= 16'h0000;
            12'd40 : o_data <= 16'h0000;
            12'd41 : o_data <= 16'h0000;
            12'd42 : o_data <= 16'h0000;
            12'd43 : o_data <= 16'h0000;
            12'd44 : o_data <= 16'h0000;
            12'd45 : o_data <= 16'h0000;
            12'd46 : o_data <= 16'h0000;
            12'd47 : o_data <= 16'h0000;
            12'd48 : o_data <= 16'h0000;
            12'd49 : o_data <= 16'h0000;
            12'd50 : o_data <= 16'h0000;
            12'd51 : o_data <= 16'h0000;
            12'd52 : o_data <= 16'h0000;
            12'd53 : o_data <= 16'h0000;
            12'd54 : o_data <= 16'h0000;
            12'd55 : o_data <= 16'h0000;
            12'd56 : o_data <= 16'h0000;
            12'd57 : o_data <= 16'h0000;
            12'd58 : o_data <= 16'h0000;
            12'd59 : o_data <= 16'h0000;
            12'd60 : o_data <= 16'h0000;
            12'd61 : o_data <= 16'h0000;
            12'd62 : o_data <= 16'h0000;
            12'd63 : o_data <= 16'h0000;
            12'd64 : o_data <= 16'h0000;
            12'd65 : o_data <= 16'h0000;
            12'd66 : o_data <= 16'h0000;
            12'd67 : o_data <= 16'h0000;
            12'd68 : o_data <= 16'h0000;
            12'd69 : o_data <= 16'h0000;
            12'd70 : o_data <= 16'h0000;
            12'd71 : o_data <= 16'h0000;
            12'd72 : o_data <= 16'h0000;
            12'd73 : o_data <= 16'h0000;
            12'd74 : o_data <= 16'h0000;
            12'd75 : o_data <= 16'h0000;
            12'd76 : o_data <= 16'h0000;
            12'd77 : o_data <= 16'h0000;
            12'd78 : o_data <= 16'h0000;
            12'd79 : o_data <= 16'h0000;
            12'd80 : o_data <= 16'h0000;
            12'd81 : o_data <= 16'h0000;
            12'd82 : o_data <= 16'h0000;
            12'd83 : o_data <= 16'h0000;
            12'd84 : o_data <= 16'h0000;
            12'd85 : o_data <= 16'h0000;
            12'd86 : o_data <= 16'h0000;
            12'd87 : o_data <= 16'h0000;
            12'd88 : o_data <= 16'h0000;
            12'd89 : o_data <= 16'h0000;
            12'd90 : o_data <= 16'h0000;
            12'd91 : o_data <= 16'h0000;
            12'd92 : o_data <= 16'h0000;
            12'd93 : o_data <= 16'h0000;
            12'd94 : o_data <= 16'h0000;
            12'd95 : o_data <= 16'h0000;
            12'd96 : o_data <= 16'h0000;
            12'd97 : o_data <= 16'h0000;
            12'd98 : o_data <= 16'h0000;
            12'd99 : o_data <= 16'h0000;
            12'd100 : o_data <= 16'h0000;
            12'd101 : o_data <= 16'h0000;
            12'd102 : o_data <= 16'h0000;
            12'd103 : o_data <= 16'h0000;
            12'd104 : o_data <= 16'h0000;
            12'd105 : o_data <= 16'h0000;
            12'd106 : o_data <= 16'h0000;
            12'd107 : o_data <= 16'h0000;
            12'd108 : o_data <= 16'h0000;
            12'd109 : o_data <= 16'h0000;
            12'd110 : o_data <= 16'h0000;
            12'd111 : o_data <= 16'h0000;
            12'd112 : o_data <= 16'h0000;
            12'd113 : o_data <= 16'h0000;
            12'd114 : o_data <= 16'h0000;
            12'd115 : o_data <= 16'h0000;
            12'd116 : o_data <= 16'h0000;
            12'd117 : o_data <= 16'h0000;
            12'd118 : o_data <= 16'h0000;
            12'd119 : o_data <= 16'h0000;
            12'd120 : o_data <= 16'h0000;
            12'd121 : o_data <= 16'h0000;
            12'd122 : o_data <= 16'h0000;
            12'd123 : o_data <= 16'h0000;
            12'd124 : o_data <= 16'h0000;
            12'd125 : o_data <= 16'h0000;
            12'd126 : o_data <= 16'h0000;
            12'd127 : o_data <= 16'h0000;
            12'd128 : o_data <= 16'h0000;
            12'd129 : o_data <= 16'h0000;
            12'd130 : o_data <= 16'h0000;
            12'd131 : o_data <= 16'h0000;
            12'd132 : o_data <= 16'h0000;
            12'd133 : o_data <= 16'h0000;
            12'd134 : o_data <= 16'h0000;
            12'd135 : o_data <= 16'h0000;
            12'd136 : o_data <= 16'h0000;
            12'd137 : o_data <= 16'h0000;
            12'd138 : o_data <= 16'h0000;
            12'd139 : o_data <= 16'h0000;
            12'd140 : o_data <= 16'h0000;
            12'd141 : o_data <= 16'h0000;
            12'd142 : o_data <= 16'h0000;
            12'd143 : o_data <= 16'h0000;
            12'd144 : o_data <= 16'h0000;
            12'd145 : o_data <= 16'h0000;
            12'd146 : o_data <= 16'h0000;
            12'd147 : o_data <= 16'h0000;
            12'd148 : o_data <= 16'h0000;
            12'd149 : o_data <= 16'h0000;
            12'd150 : o_data <= 16'h0000;
            12'd151 : o_data <= 16'h0000;
            12'd152 : o_data <= 16'h0000;
            12'd153 : o_data <= 16'h0000;
            12'd154 : o_data <= 16'h0000;
            12'd155 : o_data <= 16'h0000;
            12'd156 : o_data <= 16'h0000;
            12'd157 : o_data <= 16'h0000;
            12'd158 : o_data <= 16'h0000;
            12'd159 : o_data <= 16'h0000;
            12'd160 : o_data <= 16'h0000;
            12'd161 : o_data <= 16'h0000;
            12'd162 : o_data <= 16'h0000;
            12'd163 : o_data <= 16'h0000;
            12'd164 : o_data <= 16'h0000;
            12'd165 : o_data <= 16'h0000;
            12'd166 : o_data <= 16'h0000;
            12'd167 : o_data <= 16'h0000;
            12'd168 : o_data <= 16'h0000;
            12'd169 : o_data <= 16'h0000;
            12'd170 : o_data <= 16'h0000;
            12'd171 : o_data <= 16'h0000;
            12'd172 : o_data <= 16'h0000;
            12'd173 : o_data <= 16'h0000;
            12'd174 : o_data <= 16'h0000;
            12'd175 : o_data <= 16'h0000;
            12'd176 : o_data <= 16'h0000;
            12'd177 : o_data <= 16'h0000;
            12'd178 : o_data <= 16'h0000;
            12'd179 : o_data <= 16'h0000;
            12'd180 : o_data <= 16'h0000;
            12'd181 : o_data <= 16'h0000;
            12'd182 : o_data <= 16'h0000;
            12'd183 : o_data <= 16'h0000;
            12'd184 : o_data <= 16'h0000;
            12'd185 : o_data <= 16'h0000;
            12'd186 : o_data <= 16'h0000;
            12'd187 : o_data <= 16'h0000;
            12'd188 : o_data <= 16'h0000;
            12'd189 : o_data <= 16'h0000;
            12'd190 : o_data <= 16'h0000;
            12'd191 : o_data <= 16'h0000;
            12'd192 : o_data <= 16'h0000;
            12'd193 : o_data <= 16'h0000;
            12'd194 : o_data <= 16'h0000;
            12'd195 : o_data <= 16'h0000;
            12'd196 : o_data <= 16'h0000;
            12'd197 : o_data <= 16'h0000;
            12'd198 : o_data <= 16'h0000;
            12'd199 : o_data <= 16'h0000;
            12'd200 : o_data <= 16'h0000;
            12'd201 : o_data <= 16'h0000;
            12'd202 : o_data <= 16'h0000;
            12'd203 : o_data <= 16'h0000;
            12'd204 : o_data <= 16'h0000;
            12'd205 : o_data <= 16'h0000;
            12'd206 : o_data <= 16'h0000;
            12'd207 : o_data <= 16'h0000;
            12'd208 : o_data <= 16'h0000;
            12'd209 : o_data <= 16'h0000;
            12'd210 : o_data <= 16'h0000;
            12'd211 : o_data <= 16'h0000;
            12'd212 : o_data <= 16'h0000;
            12'd213 : o_data <= 16'h0000;
            12'd214 : o_data <= 16'h0000;
            12'd215 : o_data <= 16'h0000;
            12'd216 : o_data <= 16'h0000;
            12'd217 : o_data <= 16'h0000;
            12'd218 : o_data <= 16'h0000;
            12'd219 : o_data <= 16'h0000;
            12'd220 : o_data <= 16'h0000;
            12'd221 : o_data <= 16'h0000;
            12'd222 : o_data <= 16'h0000;
            12'd223 : o_data <= 16'h0000;
            12'd224 : o_data <= 16'h0000;
            12'd225 : o_data <= 16'h0000;
            12'd226 : o_data <= 16'h0000;
            12'd227 : o_data <= 16'h0000;
            12'd228 : o_data <= 16'h0000;
            12'd229 : o_data <= 16'h0000;
            12'd230 : o_data <= 16'h0000;
            12'd231 : o_data <= 16'h0000;
            12'd232 : o_data <= 16'h0000;
            12'd233 : o_data <= 16'h0000;
            12'd234 : o_data <= 16'h0000;
            12'd235 : o_data <= 16'h0000;
            12'd236 : o_data <= 16'h0000;
            12'd237 : o_data <= 16'h0000;
            12'd238 : o_data <= 16'h0000;
            12'd239 : o_data <= 16'h0000;
            12'd240 : o_data <= 16'h0000;
            12'd241 : o_data <= 16'h0000;
            12'd242 : o_data <= 16'h0000;
            12'd243 : o_data <= 16'h0000;
            12'd244 : o_data <= 16'h0000;
            12'd245 : o_data <= 16'h0000;
            12'd246 : o_data <= 16'h0000;
            12'd247 : o_data <= 16'h0000;
            12'd248 : o_data <= 16'h0000;
            12'd249 : o_data <= 16'h0000;
            12'd250 : o_data <= 16'h0000;
            12'd251 : o_data <= 16'h0000;
            12'd252 : o_data <= 16'h0000;
            12'd253 : o_data <= 16'h0000;
            12'd254 : o_data <= 16'h0000;
            12'd255 : o_data <= 16'h0000;
            12'd256 : o_data <= 16'h0000;
            12'd257 : o_data <= 16'h0000;
            12'd258 : o_data <= 16'h0000;
            12'd259 : o_data <= 16'h0000;
            12'd260 : o_data <= 16'h0000;
            12'd261 : o_data <= 16'h0000;
            12'd262 : o_data <= 16'h0000;
            12'd263 : o_data <= 16'h0000;
            12'd264 : o_data <= 16'h0000;
            12'd265 : o_data <= 16'h0000;
            12'd266 : o_data <= 16'h0000;
            12'd267 : o_data <= 16'h0000;
            12'd268 : o_data <= 16'h0000;
            12'd269 : o_data <= 16'h0000;
            12'd270 : o_data <= 16'h0000;
            12'd271 : o_data <= 16'h0000;
            12'd272 : o_data <= 16'h0000;
            12'd273 : o_data <= 16'h0000;
            12'd274 : o_data <= 16'h0000;
            12'd275 : o_data <= 16'h0000;
            12'd276 : o_data <= 16'h0000;
            12'd277 : o_data <= 16'h0000;
            12'd278 : o_data <= 16'h0000;
            12'd279 : o_data <= 16'h0000;
            12'd280 : o_data <= 16'h0000;
            12'd281 : o_data <= 16'h0000;
            12'd282 : o_data <= 16'h0000;
            12'd283 : o_data <= 16'h0000;
            12'd284 : o_data <= 16'h0000;
            12'd285 : o_data <= 16'h0000;
            12'd286 : o_data <= 16'h0000;
            12'd287 : o_data <= 16'h0000;
            12'd288 : o_data <= 16'h0000;
            12'd289 : o_data <= 16'h0000;
            12'd290 : o_data <= 16'h0000;
            12'd291 : o_data <= 16'h0000;
            12'd292 : o_data <= 16'h0000;
            12'd293 : o_data <= 16'h0000;
            12'd294 : o_data <= 16'h0000;
            12'd295 : o_data <= 16'h0000;
            12'd296 : o_data <= 16'h0000;
            12'd297 : o_data <= 16'h0000;
            12'd298 : o_data <= 16'h0000;
            12'd299 : o_data <= 16'h0000;
            12'd300 : o_data <= 16'h0000;
            12'd301 : o_data <= 16'h0000;
            12'd302 : o_data <= 16'h0000;
            12'd303 : o_data <= 16'h0000;
            12'd304 : o_data <= 16'h0000;
            12'd305 : o_data <= 16'h0000;
            12'd306 : o_data <= 16'h0000;
            12'd307 : o_data <= 16'h0000;
            12'd308 : o_data <= 16'h0000;
            12'd309 : o_data <= 16'h0000;
            12'd310 : o_data <= 16'h0000;
            12'd311 : o_data <= 16'h0000;
            12'd312 : o_data <= 16'h0000;
            12'd313 : o_data <= 16'h0000;
            12'd314 : o_data <= 16'h0000;
            12'd315 : o_data <= 16'h0000;
            12'd316 : o_data <= 16'h0000;
            12'd317 : o_data <= 16'h0000;
            12'd318 : o_data <= 16'h0000;
            12'd319 : o_data <= 16'h0000;
            12'd320 : o_data <= 16'h0000;
            12'd321 : o_data <= 16'h0000;
            12'd322 : o_data <= 16'h0000;
            12'd323 : o_data <= 16'h0000;
            12'd324 : o_data <= 16'h0000;
            12'd325 : o_data <= 16'h0000;
            12'd326 : o_data <= 16'h0000;
            12'd327 : o_data <= 16'h0000;
            12'd328 : o_data <= 16'h0000;
            12'd329 : o_data <= 16'h0000;
            12'd330 : o_data <= 16'h0000;
            12'd331 : o_data <= 16'h0000;
            12'd332 : o_data <= 16'h0000;
            12'd333 : o_data <= 16'h0000;
            12'd334 : o_data <= 16'h0000;
            12'd335 : o_data <= 16'h0000;
            12'd336 : o_data <= 16'h0000;
            12'd337 : o_data <= 16'h0000;
            12'd338 : o_data <= 16'h0000;
            12'd339 : o_data <= 16'h0000;
            12'd340 : o_data <= 16'h0000;
            12'd341 : o_data <= 16'h0000;
            12'd342 : o_data <= 16'h0000;
            12'd343 : o_data <= 16'h0000;
            12'd344 : o_data <= 16'h0000;
            12'd345 : o_data <= 16'h0000;
            12'd346 : o_data <= 16'h0000;
            12'd347 : o_data <= 16'h0000;
            12'd348 : o_data <= 16'h0000;
            12'd349 : o_data <= 16'h0000;
            12'd350 : o_data <= 16'h0000;
            12'd351 : o_data <= 16'h0000;
            12'd352 : o_data <= 16'h0000;
            12'd353 : o_data <= 16'h0000;
            12'd354 : o_data <= 16'h0000;
            12'd355 : o_data <= 16'h0000;
            12'd356 : o_data <= 16'h0000;
            12'd357 : o_data <= 16'h0000;
            12'd358 : o_data <= 16'h0000;
            12'd359 : o_data <= 16'h0000;
            12'd360 : o_data <= 16'h0000;
            12'd361 : o_data <= 16'h0000;
            12'd362 : o_data <= 16'h0000;
            12'd363 : o_data <= 16'h0000;
            12'd364 : o_data <= 16'h0000;
            12'd365 : o_data <= 16'h0000;
            12'd366 : o_data <= 16'h0000;
            12'd367 : o_data <= 16'h0000;
            12'd368 : o_data <= 16'h0000;
            12'd369 : o_data <= 16'h0000;
            12'd370 : o_data <= 16'h0000;
            12'd371 : o_data <= 16'h0000;
            12'd372 : o_data <= 16'h0000;
            12'd373 : o_data <= 16'h0000;
            12'd374 : o_data <= 16'h0000;
            12'd375 : o_data <= 16'h0000;
            12'd376 : o_data <= 16'h0000;
            12'd377 : o_data <= 16'h0000;
            12'd378 : o_data <= 16'h0000;
            12'd379 : o_data <= 16'h0000;
            12'd380 : o_data <= 16'h0000;
            12'd381 : o_data <= 16'h0000;
            12'd382 : o_data <= 16'h0000;
            12'd383 : o_data <= 16'h0000;
            12'd384 : o_data <= 16'h0000;
            12'd385 : o_data <= 16'h0000;
            12'd386 : o_data <= 16'h0000;
            12'd387 : o_data <= 16'h0000;
            12'd388 : o_data <= 16'h0000;
            12'd389 : o_data <= 16'h0000;
            12'd390 : o_data <= 16'h0000;
            12'd391 : o_data <= 16'h0000;
            12'd392 : o_data <= 16'h0000;
            12'd393 : o_data <= 16'h0000;
            12'd394 : o_data <= 16'h0000;
            12'd395 : o_data <= 16'h0000;
            12'd396 : o_data <= 16'h0000;
            12'd397 : o_data <= 16'h0000;
            12'd398 : o_data <= 16'h0000;
            12'd399 : o_data <= 16'h0000;
            12'd400 : o_data <= 16'h0000;
            12'd401 : o_data <= 16'h0000;
            12'd402 : o_data <= 16'h1860;
            12'd403 : o_data <= 16'h69C5;
            12'd404 : o_data <= 16'h7A46;
            12'd405 : o_data <= 16'h82C8;
            12'd406 : o_data <= 16'h7B2B;
            12'd407 : o_data <= 16'h838C;
            12'd408 : o_data <= 16'h7BAE;
            12'd409 : o_data <= 16'h83AE;
            12'd410 : o_data <= 16'h7B2C;
            12'd411 : o_data <= 16'h5A07;
            12'd412 : o_data <= 16'h0821;
            12'd413 : o_data <= 16'h0000;
            12'd414 : o_data <= 16'h0000;
            12'd415 : o_data <= 16'h0000;
            12'd416 : o_data <= 16'h0000;
            12'd417 : o_data <= 16'h0000;
            12'd418 : o_data <= 16'h0000;
            12'd419 : o_data <= 16'h0000;
            12'd420 : o_data <= 16'h0000;
            12'd421 : o_data <= 16'h0000;
            12'd422 : o_data <= 16'h0000;
            12'd423 : o_data <= 16'h0000;
            12'd424 : o_data <= 16'h0000;
            12'd425 : o_data <= 16'h0000;
            12'd426 : o_data <= 16'h0000;
            12'd427 : o_data <= 16'h0000;
            12'd428 : o_data <= 16'h0000;
            12'd429 : o_data <= 16'h0000;
            12'd430 : o_data <= 16'h0000;
            12'd431 : o_data <= 16'h0000;
            12'd432 : o_data <= 16'h0000;
            12'd433 : o_data <= 16'h0000;
            12'd434 : o_data <= 16'h0000;
            12'd435 : o_data <= 16'h0000;
            12'd436 : o_data <= 16'h0000;
            12'd437 : o_data <= 16'h0000;
            12'd438 : o_data <= 16'h0000;
            12'd439 : o_data <= 16'h0000;
            12'd440 : o_data <= 16'h0000;
            12'd441 : o_data <= 16'h0000;
            12'd442 : o_data <= 16'h0000;
            12'd443 : o_data <= 16'h0000;
            12'd444 : o_data <= 16'h0000;
            12'd445 : o_data <= 16'h0000;
            12'd446 : o_data <= 16'h5143;
            12'd447 : o_data <= 16'hAB88;
            12'd448 : o_data <= 16'hFD2E;
            12'd449 : o_data <= 16'hFDD0;
            12'd450 : o_data <= 16'hFDF0;
            12'd451 : o_data <= 16'hFDF1;
            12'd452 : o_data <= 16'hFE32;
            12'd453 : o_data <= 16'hFEB5;
            12'd454 : o_data <= 16'hFF16;
            12'd455 : o_data <= 16'hFEF7;
            12'd456 : o_data <= 16'hFEF6;
            12'd457 : o_data <= 16'hFEF6;
            12'd458 : o_data <= 16'hFED5;
            12'd459 : o_data <= 16'hFED5;
            12'd460 : o_data <= 16'hFF17;
            12'd461 : o_data <= 16'hFED6;
            12'd462 : o_data <= 16'hE551;
            12'd463 : o_data <= 16'h934A;
            12'd464 : o_data <= 16'h5165;
            12'd465 : o_data <= 16'h0000;
            12'd466 : o_data <= 16'h0000;
            12'd467 : o_data <= 16'h0000;
            12'd468 : o_data <= 16'h0000;
            12'd469 : o_data <= 16'h0000;
            12'd470 : o_data <= 16'h0000;
            12'd471 : o_data <= 16'h0000;
            12'd472 : o_data <= 16'h0000;
            12'd473 : o_data <= 16'h0000;
            12'd474 : o_data <= 16'h0000;
            12'd475 : o_data <= 16'h0000;
            12'd476 : o_data <= 16'h0000;
            12'd477 : o_data <= 16'h0000;
            12'd478 : o_data <= 16'h0000;
            12'd479 : o_data <= 16'h0000;
            12'd480 : o_data <= 16'h0000;
            12'd481 : o_data <= 16'h0000;
            12'd482 : o_data <= 16'h0000;
            12'd483 : o_data <= 16'h0000;
            12'd484 : o_data <= 16'h0000;
            12'd485 : o_data <= 16'h0000;
            12'd486 : o_data <= 16'h0000;
            12'd487 : o_data <= 16'h0000;
            12'd488 : o_data <= 16'h0000;
            12'd489 : o_data <= 16'h0000;
            12'd490 : o_data <= 16'h0000;
            12'd491 : o_data <= 16'h0000;
            12'd492 : o_data <= 16'h7A65;
            12'd493 : o_data <= 16'hFDB0;
            12'd494 : o_data <= 16'hFE52;
            12'd495 : o_data <= 16'hFDD2;
            12'd496 : o_data <= 16'hFD92;
            12'd497 : o_data <= 16'hFD71;
            12'd498 : o_data <= 16'hFD30;
            12'd499 : o_data <= 16'hF590;
            12'd500 : o_data <= 16'hFDB1;
            12'd501 : o_data <= 16'hFD4E;
            12'd502 : o_data <= 16'hF52D;
            12'd503 : o_data <= 16'hFD6D;
            12'd504 : o_data <= 16'hFD8E;
            12'd505 : o_data <= 16'hF5AE;
            12'd506 : o_data <= 16'hFDCF;
            12'd507 : o_data <= 16'hF5F0;
            12'd508 : o_data <= 16'hF5F0;
            12'd509 : o_data <= 16'hF5D1;
            12'd510 : o_data <= 16'hFDF1;
            12'd511 : o_data <= 16'hFDF1;
            12'd512 : o_data <= 16'hFE12;
            12'd513 : o_data <= 16'hFE32;
            12'd514 : o_data <= 16'hCC2C;
            12'd515 : o_data <= 16'h5143;
            12'd516 : o_data <= 16'h0000;
            12'd517 : o_data <= 16'h0000;
            12'd518 : o_data <= 16'h0000;
            12'd519 : o_data <= 16'h0000;
            12'd520 : o_data <= 16'h0000;
            12'd521 : o_data <= 16'h0000;
            12'd522 : o_data <= 16'h0000;
            12'd523 : o_data <= 16'h0000;
            12'd524 : o_data <= 16'h0000;
            12'd525 : o_data <= 16'h0000;
            12'd526 : o_data <= 16'h0000;
            12'd527 : o_data <= 16'h0000;
            12'd528 : o_data <= 16'h0000;
            12'd529 : o_data <= 16'h0000;
            12'd530 : o_data <= 16'h0000;
            12'd531 : o_data <= 16'h0000;
            12'd532 : o_data <= 16'h0000;
            12'd533 : o_data <= 16'h0000;
            12'd534 : o_data <= 16'h0000;
            12'd535 : o_data <= 16'h0000;
            12'd536 : o_data <= 16'h0000;
            12'd537 : o_data <= 16'h0000;
            12'd538 : o_data <= 16'h0000;
            12'd539 : o_data <= 16'hFD6F;
            12'd540 : o_data <= 16'hFE74;
            12'd541 : o_data <= 16'hFD91;
            12'd542 : o_data <= 16'hFC8D;
            12'd543 : o_data <= 16'hFC2B;
            12'd544 : o_data <= 16'hFC4A;
            12'd545 : o_data <= 16'hF429;
            12'd546 : o_data <= 16'hFD0C;
            12'd547 : o_data <= 16'hF4CA;
            12'd548 : o_data <= 16'hFC88;
            12'd549 : o_data <= 16'hF4A9;
            12'd550 : o_data <= 16'hFCC9;
            12'd551 : o_data <= 16'hF4E9;
            12'd552 : o_data <= 16'hFD08;
            12'd553 : o_data <= 16'hFD09;
            12'd554 : o_data <= 16'hF509;
            12'd555 : o_data <= 16'hFD09;
            12'd556 : o_data <= 16'hF509;
            12'd557 : o_data <= 16'hFD2B;
            12'd558 : o_data <= 16'hF5AE;
            12'd559 : o_data <= 16'hF5AE;
            12'd560 : o_data <= 16'hF5B0;
            12'd561 : o_data <= 16'hF5D1;
            12'd562 : o_data <= 16'hFDF2;
            12'd563 : o_data <= 16'hFE12;
            12'd564 : o_data <= 16'hFCEE;
            12'd565 : o_data <= 16'h5143;
            12'd566 : o_data <= 16'h0000;
            12'd567 : o_data <= 16'h0000;
            12'd568 : o_data <= 16'h0000;
            12'd569 : o_data <= 16'h0000;
            12'd570 : o_data <= 16'h0000;
            12'd571 : o_data <= 16'h0000;
            12'd572 : o_data <= 16'h0000;
            12'd573 : o_data <= 16'h0000;
            12'd574 : o_data <= 16'h0000;
            12'd575 : o_data <= 16'h0000;
            12'd576 : o_data <= 16'h0000;
            12'd577 : o_data <= 16'h0000;
            12'd578 : o_data <= 16'h0000;
            12'd579 : o_data <= 16'h0000;
            12'd580 : o_data <= 16'h0000;
            12'd581 : o_data <= 16'h0000;
            12'd582 : o_data <= 16'h0000;
            12'd583 : o_data <= 16'h0000;
            12'd584 : o_data <= 16'h0000;
            12'd585 : o_data <= 16'h1840;
            12'd586 : o_data <= 16'hFEB3;
            12'd587 : o_data <= 16'hFE54;
            12'd588 : o_data <= 16'hFC8D;
            12'd589 : o_data <= 16'hFC4A;
            12'd590 : o_data <= 16'hFC89;
            12'd591 : o_data <= 16'hFC88;
            12'd592 : o_data <= 16'hFC86;
            12'd593 : o_data <= 16'hFDAD;
            12'd594 : o_data <= 16'hF528;
            12'd595 : o_data <= 16'hFD07;
            12'd596 : o_data <= 16'hFD27;
            12'd597 : o_data <= 16'hFD27;
            12'd598 : o_data <= 16'hFD47;
            12'd599 : o_data <= 16'hFD27;
            12'd600 : o_data <= 16'hF507;
            12'd601 : o_data <= 16'hFD07;
            12'd602 : o_data <= 16'hFCC6;
            12'd603 : o_data <= 16'hF54B;
            12'd604 : o_data <= 16'hFDAC;
            12'd605 : o_data <= 16'hF52A;
            12'd606 : o_data <= 16'hF4A7;
            12'd607 : o_data <= 16'hFCA8;
            12'd608 : o_data <= 16'hF4A8;
            12'd609 : o_data <= 16'hF4AA;
            12'd610 : o_data <= 16'hF50C;
            12'd611 : o_data <= 16'hF54E;
            12'd612 : o_data <= 16'hFDB1;
            12'd613 : o_data <= 16'hFDB0;
            12'd614 : o_data <= 16'hE40A;
            12'd615 : o_data <= 16'h0000;
            12'd616 : o_data <= 16'h0000;
            12'd617 : o_data <= 16'h0000;
            12'd618 : o_data <= 16'h0000;
            12'd619 : o_data <= 16'h0000;
            12'd620 : o_data <= 16'h0000;
            12'd621 : o_data <= 16'h0000;
            12'd622 : o_data <= 16'h0000;
            12'd623 : o_data <= 16'h0000;
            12'd624 : o_data <= 16'h0000;
            12'd625 : o_data <= 16'h0000;
            12'd626 : o_data <= 16'h0000;
            12'd627 : o_data <= 16'h0000;
            12'd628 : o_data <= 16'h0000;
            12'd629 : o_data <= 16'h0000;
            12'd630 : o_data <= 16'h0000;
            12'd631 : o_data <= 16'h0000;
            12'd632 : o_data <= 16'h0000;
            12'd633 : o_data <= 16'hFE72;
            12'd634 : o_data <= 16'hFDF3;
            12'd635 : o_data <= 16'hFCA9;
            12'd636 : o_data <= 16'hFD08;
            12'd637 : o_data <= 16'hFD48;
            12'd638 : o_data <= 16'hFD66;
            12'd639 : o_data <= 16'hFE2B;
            12'd640 : o_data <= 16'hF60C;
            12'd641 : o_data <= 16'hFD46;
            12'd642 : o_data <= 16'hFD05;
            12'd643 : o_data <= 16'hFCE5;
            12'd644 : o_data <= 16'hFD05;
            12'd645 : o_data <= 16'hFCE5;
            12'd646 : o_data <= 16'hF4C5;
            12'd647 : o_data <= 16'hFD87;
            12'd648 : o_data <= 16'hFE4B;
            12'd649 : o_data <= 16'hF6B0;
            12'd650 : o_data <= 16'hFEAF;
            12'd651 : o_data <= 16'hFDC8;
            12'd652 : o_data <= 16'hFD26;
            12'd653 : o_data <= 16'hFCE7;
            12'd654 : o_data <= 16'hFCC7;
            12'd655 : o_data <= 16'hF4A8;
            12'd656 : o_data <= 16'hFC87;
            12'd657 : o_data <= 16'hF487;
            12'd658 : o_data <= 16'hFC68;
            12'd659 : o_data <= 16'hF489;
            12'd660 : o_data <= 16'hF4CB;
            12'd661 : o_data <= 16'hF56F;
            12'd662 : o_data <= 16'hFD70;
            12'd663 : o_data <= 16'hFD8E;
            12'd664 : o_data <= 16'h28C2;
            12'd665 : o_data <= 16'h0000;
            12'd666 : o_data <= 16'h0000;
            12'd667 : o_data <= 16'h0000;
            12'd668 : o_data <= 16'h0000;
            12'd669 : o_data <= 16'h0000;
            12'd670 : o_data <= 16'h0000;
            12'd671 : o_data <= 16'h0000;
            12'd672 : o_data <= 16'h0000;
            12'd673 : o_data <= 16'h0000;
            12'd674 : o_data <= 16'h0000;
            12'd675 : o_data <= 16'h0000;
            12'd676 : o_data <= 16'h0000;
            12'd677 : o_data <= 16'h0000;
            12'd678 : o_data <= 16'h0000;
            12'd679 : o_data <= 16'h0000;
            12'd680 : o_data <= 16'h9B48;
            12'd681 : o_data <= 16'hFEB4;
            12'd682 : o_data <= 16'hFD68;
            12'd683 : o_data <= 16'hFDA8;
            12'd684 : o_data <= 16'hFD86;
            12'd685 : o_data <= 16'hFCA5;
            12'd686 : o_data <= 16'hFD09;
            12'd687 : o_data <= 16'hFB43;
            12'd688 : o_data <= 16'hFAE3;
            12'd689 : o_data <= 16'hFAA3;
            12'd690 : o_data <= 16'hFA62;
            12'd691 : o_data <= 16'hFA42;
            12'd692 : o_data <= 16'hFA62;
            12'd693 : o_data <= 16'hFB24;
            12'd694 : o_data <= 16'hFB86;
            12'd695 : o_data <= 16'hFAE3;
            12'd696 : o_data <= 16'hFAC1;
            12'd697 : o_data <= 16'hFAA0;
            12'd698 : o_data <= 16'hFB61;
            12'd699 : o_data <= 16'hFC85;
            12'd700 : o_data <= 16'hF5A8;
            12'd701 : o_data <= 16'hFE09;
            12'd702 : o_data <= 16'hFD87;
            12'd703 : o_data <= 16'hFD07;
            12'd704 : o_data <= 16'hF4C6;
            12'd705 : o_data <= 16'hFC87;
            12'd706 : o_data <= 16'hF467;
            12'd707 : o_data <= 16'hFC67;
            12'd708 : o_data <= 16'hFC48;
            12'd709 : o_data <= 16'hFC6A;
            12'd710 : o_data <= 16'hF4EC;
            12'd711 : o_data <= 16'hFD4F;
            12'd712 : o_data <= 16'hFDAF;
            12'd713 : o_data <= 16'h69A3;
            12'd714 : o_data <= 16'h0000;
            12'd715 : o_data <= 16'h0000;
            12'd716 : o_data <= 16'h0000;
            12'd717 : o_data <= 16'h0000;
            12'd718 : o_data <= 16'h0000;
            12'd719 : o_data <= 16'h0000;
            12'd720 : o_data <= 16'h0000;
            12'd721 : o_data <= 16'h0000;
            12'd722 : o_data <= 16'h0000;
            12'd723 : o_data <= 16'h0000;
            12'd724 : o_data <= 16'h0000;
            12'd725 : o_data <= 16'h0000;
            12'd726 : o_data <= 16'h0000;
            12'd727 : o_data <= 16'h0000;
            12'd728 : o_data <= 16'hFF17;
            12'd729 : o_data <= 16'hFD46;
            12'd730 : o_data <= 16'hFCC5;
            12'd731 : o_data <= 16'hFB84;
            12'd732 : o_data <= 16'hFAC3;
            12'd733 : o_data <= 16'hFBC7;
            12'd734 : o_data <= 16'hF9C1;
            12'd735 : o_data <= 16'hF9A1;
            12'd736 : o_data <= 16'hF960;
            12'd737 : o_data <= 16'hF100;
            12'd738 : o_data <= 16'hE8E0;
            12'd739 : o_data <= 16'hF9E2;
            12'd740 : o_data <= 16'hE9A2;
            12'd741 : o_data <= 16'hF100;
            12'd742 : o_data <= 16'hF120;
            12'd743 : o_data <= 16'hE961;
            12'd744 : o_data <= 16'hF1A1;
            12'd745 : o_data <= 16'hFA02;
            12'd746 : o_data <= 16'hFA01;
            12'd747 : o_data <= 16'hFA01;
            12'd748 : o_data <= 16'hFA60;
            12'd749 : o_data <= 16'hFB41;
            12'd750 : o_data <= 16'hFCE5;
            12'd751 : o_data <= 16'hFE0B;
            12'd752 : o_data <= 16'hFDEB;
            12'd753 : o_data <= 16'hFD69;
            12'd754 : o_data <= 16'hFD29;
            12'd755 : o_data <= 16'hF50A;
            12'd756 : o_data <= 16'hF50B;
            12'd757 : o_data <= 16'hFD0C;
            12'd758 : o_data <= 16'hF56E;
            12'd759 : o_data <= 16'hFD2F;
            12'd760 : o_data <= 16'hF54F;
            12'd761 : o_data <= 16'hFDCF;
            12'd762 : o_data <= 16'h30C2;
            12'd763 : o_data <= 16'h0000;
            12'd764 : o_data <= 16'h0000;
            12'd765 : o_data <= 16'h0000;
            12'd766 : o_data <= 16'h0000;
            12'd767 : o_data <= 16'h0000;
            12'd768 : o_data <= 16'h0000;
            12'd769 : o_data <= 16'h0000;
            12'd770 : o_data <= 16'h0000;
            12'd771 : o_data <= 16'h0000;
            12'd772 : o_data <= 16'h0000;
            12'd773 : o_data <= 16'h0000;
            12'd774 : o_data <= 16'h0000;
            12'd775 : o_data <= 16'h1841;
            12'd776 : o_data <= 16'hFD09;
            12'd777 : o_data <= 16'hFB23;
            12'd778 : o_data <= 16'hFA42;
            12'd779 : o_data <= 16'hF940;
            12'd780 : o_data <= 16'hFA42;
            12'd781 : o_data <= 16'hD101;
            12'd782 : o_data <= 16'hBA05;
            12'd783 : o_data <= 16'hAAE9;
            12'd784 : o_data <= 16'hABED;
            12'd785 : o_data <= 16'h93ED;
            12'd786 : o_data <= 16'h9C6F;
            12'd787 : o_data <= 16'h9CD1;
            12'd788 : o_data <= 16'hAD53;
            12'd789 : o_data <= 16'h9CF2;
            12'd790 : o_data <= 16'hACB1;
            12'd791 : o_data <= 16'hA40E;
            12'd792 : o_data <= 16'hB36D;
            12'd793 : o_data <= 16'hB288;
            12'd794 : o_data <= 16'hC902;
            12'd795 : o_data <= 16'hD8A0;
            12'd796 : o_data <= 16'hF161;
            12'd797 : o_data <= 16'hF263;
            12'd798 : o_data <= 16'hFB06;
            12'd799 : o_data <= 16'hFB22;
            12'd800 : o_data <= 16'hFCE4;
            12'd801 : o_data <= 16'hF608;
            12'd802 : o_data <= 16'hFD88;
            12'd803 : o_data <= 16'hFD06;
            12'd804 : o_data <= 16'hFCC8;
            12'd805 : o_data <= 16'hFCA9;
            12'd806 : o_data <= 16'hFC89;
            12'd807 : o_data <= 16'hF48B;
            12'd808 : o_data <= 16'hFCED;
            12'd809 : o_data <= 16'hFD6F;
            12'd810 : o_data <= 16'hFDAF;
            12'd811 : o_data <= 16'h0000;
            12'd812 : o_data <= 16'h0000;
            12'd813 : o_data <= 16'h0000;
            12'd814 : o_data <= 16'h0000;
            12'd815 : o_data <= 16'h0000;
            12'd816 : o_data <= 16'h0000;
            12'd817 : o_data <= 16'h0000;
            12'd818 : o_data <= 16'h0000;
            12'd819 : o_data <= 16'h0000;
            12'd820 : o_data <= 16'h0000;
            12'd821 : o_data <= 16'h0000;
            12'd822 : o_data <= 16'h0000;
            12'd823 : o_data <= 16'h0000;
            12'd824 : o_data <= 16'hDA85;
            12'd825 : o_data <= 16'hE9C3;
            12'd826 : o_data <= 16'hC3AC;
            12'd827 : o_data <= 16'hB533;
            12'd828 : o_data <= 16'hBE57;
            12'd829 : o_data <= 16'hDFBD;
            12'd830 : o_data <= 16'hE77D;
            12'd831 : o_data <= 16'hC677;
            12'd832 : o_data <= 16'hDEFA;
            12'd833 : o_data <= 16'hD698;
            12'd834 : o_data <= 16'hE71B;
            12'd835 : o_data <= 16'hE6F9;
            12'd836 : o_data <= 16'hF77D;
            12'd837 : o_data <= 16'hE73B;
            12'd838 : o_data <= 16'hEF3B;
            12'd839 : o_data <= 16'hEF7D;
            12'd840 : o_data <= 16'hE71A;
            12'd841 : o_data <= 16'hD71A;
            12'd842 : o_data <= 16'hDF3B;
            12'd843 : o_data <= 16'hB594;
            12'd844 : o_data <= 16'hCCAF;
            12'd845 : o_data <= 16'hC102;
            12'd846 : o_data <= 16'hE060;
            12'd847 : o_data <= 16'hE940;
            12'd848 : o_data <= 16'hF9E2;
            12'd849 : o_data <= 16'hFB42;
            12'd850 : o_data <= 16'hFD86;
            12'd851 : o_data <= 16'hFE2A;
            12'd852 : o_data <= 16'hFD68;
            12'd853 : o_data <= 16'hFD29;
            12'd854 : o_data <= 16'hFD0A;
            12'd855 : o_data <= 16'hFCCB;
            12'd856 : o_data <= 16'hFCCC;
            12'd857 : o_data <= 16'hFD0E;
            12'd858 : o_data <= 16'hFE52;
            12'd859 : o_data <= 16'h3103;
            12'd860 : o_data <= 16'h0000;
            12'd861 : o_data <= 16'h0000;
            12'd862 : o_data <= 16'h0000;
            12'd863 : o_data <= 16'h0000;
            12'd864 : o_data <= 16'h0000;
            12'd865 : o_data <= 16'h0000;
            12'd866 : o_data <= 16'h0000;
            12'd867 : o_data <= 16'h0000;
            12'd868 : o_data <= 16'h0000;
            12'd869 : o_data <= 16'h0000;
            12'd870 : o_data <= 16'h0000;
            12'd871 : o_data <= 16'h0000;
            12'd872 : o_data <= 16'h3A8A;
            12'd873 : o_data <= 16'hD79B;
            12'd874 : o_data <= 16'hBE36;
            12'd875 : o_data <= 16'hEF9D;
            12'd876 : o_data <= 16'hE71A;
            12'd877 : o_data <= 16'hEF3C;
            12'd878 : o_data <= 16'hE71A;
            12'd879 : o_data <= 16'hEF3C;
            12'd880 : o_data <= 16'hE71A;
            12'd881 : o_data <= 16'hD6B9;
            12'd882 : o_data <= 16'hD678;
            12'd883 : o_data <= 16'hE73B;
            12'd884 : o_data <= 16'hDED9;
            12'd885 : o_data <= 16'hE71B;
            12'd886 : o_data <= 16'hE71A;
            12'd887 : o_data <= 16'hE6FA;
            12'd888 : o_data <= 16'hDEDA;
            12'd889 : o_data <= 16'hE71B;
            12'd890 : o_data <= 16'hE6FA;
            12'd891 : o_data <= 16'hE71B;
            12'd892 : o_data <= 16'hE73B;
            12'd893 : o_data <= 16'hCED9;
            12'd894 : o_data <= 16'hB553;
            12'd895 : o_data <= 16'hBA87;
            12'd896 : o_data <= 16'hE0A0;
            12'd897 : o_data <= 16'hF181;
            12'd898 : o_data <= 16'hF9C1;
            12'd899 : o_data <= 16'hFBE3;
            12'd900 : o_data <= 16'hFEAC;
            12'd901 : o_data <= 16'hFE4E;
            12'd902 : o_data <= 16'hFDEC;
            12'd903 : o_data <= 16'hFDAD;
            12'd904 : o_data <= 16'hFD6D;
            12'd905 : o_data <= 16'hFD4E;
            12'd906 : o_data <= 16'hFED4;
            12'd907 : o_data <= 16'h2924;
            12'd908 : o_data <= 16'h0000;
            12'd909 : o_data <= 16'h0000;
            12'd910 : o_data <= 16'h0000;
            12'd911 : o_data <= 16'h0000;
            12'd912 : o_data <= 16'h0000;
            12'd913 : o_data <= 16'h0000;
            12'd914 : o_data <= 16'h0000;
            12'd915 : o_data <= 16'h0000;
            12'd916 : o_data <= 16'h0000;
            12'd917 : o_data <= 16'h0000;
            12'd918 : o_data <= 16'h0000;
            12'd919 : o_data <= 16'h0000;
            12'd920 : o_data <= 16'h0000;
            12'd921 : o_data <= 16'hAD54;
            12'd922 : o_data <= 16'hD6D8;
            12'd923 : o_data <= 16'hCE36;
            12'd924 : o_data <= 16'hE73B;
            12'd925 : o_data <= 16'hBE36;
            12'd926 : o_data <= 16'hD6D9;
            12'd927 : o_data <= 16'hD71A;
            12'd928 : o_data <= 16'hCED9;
            12'd929 : o_data <= 16'hDF3B;
            12'd930 : o_data <= 16'hD6D9;
            12'd931 : o_data <= 16'hDED9;
            12'd932 : o_data <= 16'hCE97;
            12'd933 : o_data <= 16'hD6D9;
            12'd934 : o_data <= 16'hD6D9;
            12'd935 : o_data <= 16'hD6B8;
            12'd936 : o_data <= 16'hDF3A;
            12'd937 : o_data <= 16'hDEFA;
            12'd938 : o_data <= 16'hDED9;
            12'd939 : o_data <= 16'hE6FA;
            12'd940 : o_data <= 16'hE6FA;
            12'd941 : o_data <= 16'hEF3B;
            12'd942 : o_data <= 16'hEF5B;
            12'd943 : o_data <= 16'hDF1B;
            12'd944 : o_data <= 16'h9511;
            12'd945 : o_data <= 16'hB1C5;
            12'd946 : o_data <= 16'hF1C2;
            12'd947 : o_data <= 16'hF223;
            12'd948 : o_data <= 16'hFA61;
            12'd949 : o_data <= 16'hFCE4;
            12'd950 : o_data <= 16'hFDE7;
            12'd951 : o_data <= 16'hFD8A;
            12'd952 : o_data <= 16'hFD6B;
            12'd953 : o_data <= 16'hFDAE;
            12'd954 : o_data <= 16'hFE90;
            12'd955 : o_data <= 16'h0000;
            12'd956 : o_data <= 16'h0000;
            12'd957 : o_data <= 16'h0000;
            12'd958 : o_data <= 16'h0000;
            12'd959 : o_data <= 16'h0000;
            12'd960 : o_data <= 16'h0000;
            12'd961 : o_data <= 16'h0000;
            12'd962 : o_data <= 16'h0000;
            12'd963 : o_data <= 16'h0000;
            12'd964 : o_data <= 16'h0000;
            12'd965 : o_data <= 16'h0000;
            12'd966 : o_data <= 16'h0000;
            12'd967 : o_data <= 16'h0000;
            12'd968 : o_data <= 16'h0000;
            12'd969 : o_data <= 16'h0000;
            12'd970 : o_data <= 16'h4227;
            12'd971 : o_data <= 16'h9D53;
            12'd972 : o_data <= 16'hADB4;
            12'd973 : o_data <= 16'hE699;
            12'd974 : o_data <= 16'hF679;
            12'd975 : o_data <= 16'hFDD6;
            12'd976 : o_data <= 16'hFD96;
            12'd977 : o_data <= 16'hFD55;
            12'd978 : o_data <= 16'hFD34;
            12'd979 : o_data <= 16'hFD34;
            12'd980 : o_data <= 16'hFD14;
            12'd981 : o_data <= 16'hFD14;
            12'd982 : o_data <= 16'hF514;
            12'd983 : o_data <= 16'hFDB6;
            12'd984 : o_data <= 16'hF618;
            12'd985 : o_data <= 16'hF658;
            12'd986 : o_data <= 16'hE698;
            12'd987 : o_data <= 16'hDEB9;
            12'd988 : o_data <= 16'hCEF9;
            12'd989 : o_data <= 16'hD6DA;
            12'd990 : o_data <= 16'hDEFA;
            12'd991 : o_data <= 16'hDEB9;
            12'd992 : o_data <= 16'hEF3B;
            12'd993 : o_data <= 16'hC698;
            12'd994 : o_data <= 16'h9C4E;
            12'd995 : o_data <= 16'hC880;
            12'd996 : o_data <= 16'hF141;
            12'd997 : o_data <= 16'hF161;
            12'd998 : o_data <= 16'hFB23;
            12'd999 : o_data <= 16'hFD65;
            12'd1000 : o_data <= 16'hFDA8;
            12'd1001 : o_data <= 16'hFD27;
            12'd1002 : o_data <= 16'hAB08;
            12'd1003 : o_data <= 16'h0000;
            12'd1004 : o_data <= 16'h0000;
            12'd1005 : o_data <= 16'h0000;
            12'd1006 : o_data <= 16'h0000;
            12'd1007 : o_data <= 16'h0000;
            12'd1008 : o_data <= 16'h0000;
            12'd1009 : o_data <= 16'h0000;
            12'd1010 : o_data <= 16'h0000;
            12'd1011 : o_data <= 16'h0000;
            12'd1012 : o_data <= 16'h0000;
            12'd1013 : o_data <= 16'h0000;
            12'd1014 : o_data <= 16'h0000;
            12'd1015 : o_data <= 16'h0000;
            12'd1016 : o_data <= 16'h0000;
            12'd1017 : o_data <= 16'h0000;
            12'd1018 : o_data <= 16'h41C7;
            12'd1019 : o_data <= 16'hD514;
            12'd1020 : o_data <= 16'hFDF7;
            12'd1021 : o_data <= 16'hFD14;
            12'd1022 : o_data <= 16'hFCB2;
            12'd1023 : o_data <= 16'hF472;
            12'd1024 : o_data <= 16'hF430;
            12'd1025 : o_data <= 16'hF3CF;
            12'd1026 : o_data <= 16'hF38E;
            12'd1027 : o_data <= 16'hF30C;
            12'd1028 : o_data <= 16'hEB6E;
            12'd1029 : o_data <= 16'hF411;
            12'd1030 : o_data <= 16'hEBAE;
            12'd1031 : o_data <= 16'hF34E;
            12'd1032 : o_data <= 16'hEB4D;
            12'd1033 : o_data <= 16'hEB8E;
            12'd1034 : o_data <= 16'hF410;
            12'd1035 : o_data <= 16'hF4B3;
            12'd1036 : o_data <= 16'hFD75;
            12'd1037 : o_data <= 16'hFE38;
            12'd1038 : o_data <= 16'hE6B9;
            12'd1039 : o_data <= 16'hD6F9;
            12'd1040 : o_data <= 16'hD6B9;
            12'd1041 : o_data <= 16'hCE57;
            12'd1042 : o_data <= 16'hF79D;
            12'd1043 : o_data <= 16'hBE77;
            12'd1044 : o_data <= 16'h9A47;
            12'd1045 : o_data <= 16'hC8A0;
            12'd1046 : o_data <= 16'hE8A0;
            12'd1047 : o_data <= 16'hF120;
            12'd1048 : o_data <= 16'hEA60;
            12'd1049 : o_data <= 16'hD369;
            12'd1050 : o_data <= 16'h0001;
            12'd1051 : o_data <= 16'h0000;
            12'd1052 : o_data <= 16'h0000;
            12'd1053 : o_data <= 16'h0000;
            12'd1054 : o_data <= 16'h0000;
            12'd1055 : o_data <= 16'h0000;
            12'd1056 : o_data <= 16'h0000;
            12'd1057 : o_data <= 16'h0000;
            12'd1058 : o_data <= 16'h0000;
            12'd1059 : o_data <= 16'h0000;
            12'd1060 : o_data <= 16'h0000;
            12'd1061 : o_data <= 16'h0000;
            12'd1062 : o_data <= 16'h0000;
            12'd1063 : o_data <= 16'h0000;
            12'd1064 : o_data <= 16'h0000;
            12'd1065 : o_data <= 16'hF5D7;
            12'd1066 : o_data <= 16'hFE38;
            12'd1067 : o_data <= 16'hFD34;
            12'd1068 : o_data <= 16'hF451;
            12'd1069 : o_data <= 16'hF451;
            12'd1070 : o_data <= 16'hEC31;
            12'd1071 : o_data <= 16'hEC11;
            12'd1072 : o_data <= 16'hF3CF;
            12'd1073 : o_data <= 16'hEC11;
            12'd1074 : o_data <= 16'hF4B3;
            12'd1075 : o_data <= 16'hF493;
            12'd1076 : o_data <= 16'hF3CF;
            12'd1077 : o_data <= 16'hF2AB;
            12'd1078 : o_data <= 16'hF2CC;
            12'd1079 : o_data <= 16'hEACC;
            12'd1080 : o_data <= 16'hF2AB;
            12'd1081 : o_data <= 16'hF2AC;
            12'd1082 : o_data <= 16'hEA8B;
            12'd1083 : o_data <= 16'hEB2D;
            12'd1084 : o_data <= 16'hF430;
            12'd1085 : o_data <= 16'hEC72;
            12'd1086 : o_data <= 16'hFD55;
            12'd1087 : o_data <= 16'hFDF7;
            12'd1088 : o_data <= 16'hEE57;
            12'd1089 : o_data <= 16'hD697;
            12'd1090 : o_data <= 16'hCED9;
            12'd1091 : o_data <= 16'hE71B;
            12'd1092 : o_data <= 16'hDF3A;
            12'd1093 : o_data <= 16'hCEFA;
            12'd1094 : o_data <= 16'hB552;
            12'd1095 : o_data <= 16'hC5D5;
            12'd1096 : o_data <= 16'hCEFB;
            12'd1097 : o_data <= 16'hA5B5;
            12'd1098 : o_data <= 16'h0000;
            12'd1099 : o_data <= 16'h0000;
            12'd1100 : o_data <= 16'h0000;
            12'd1101 : o_data <= 16'h0000;
            12'd1102 : o_data <= 16'h0000;
            12'd1103 : o_data <= 16'h0000;
            12'd1104 : o_data <= 16'h0000;
            12'd1105 : o_data <= 16'h0000;
            12'd1106 : o_data <= 16'h0000;
            12'd1107 : o_data <= 16'h0000;
            12'd1108 : o_data <= 16'h0000;
            12'd1109 : o_data <= 16'h0000;
            12'd1110 : o_data <= 16'h0000;
            12'd1111 : o_data <= 16'h2945;
            12'd1112 : o_data <= 16'hFE9A;
            12'd1113 : o_data <= 16'hFCD3;
            12'd1114 : o_data <= 16'hF471;
            12'd1115 : o_data <= 16'hF3D0;
            12'd1116 : o_data <= 16'hEBAF;
            12'd1117 : o_data <= 16'hEBF0;
            12'd1118 : o_data <= 16'hEC51;
            12'd1119 : o_data <= 16'hEC52;
            12'd1120 : o_data <= 16'hF431;
            12'd1121 : o_data <= 16'hEB6E;
            12'd1122 : o_data <= 16'hEA6A;
            12'd1123 : o_data <= 16'hEAAB;
            12'd1124 : o_data <= 16'hEAAC;
            12'd1125 : o_data <= 16'hEACC;
            12'd1126 : o_data <= 16'hF2CB;
            12'd1127 : o_data <= 16'hEACC;
            12'd1128 : o_data <= 16'hF2AB;
            12'd1129 : o_data <= 16'hF3AF;
            12'd1130 : o_data <= 16'hF411;
            12'd1131 : o_data <= 16'hF3AF;
            12'd1132 : o_data <= 16'hEAAB;
            12'd1133 : o_data <= 16'hF2EC;
            12'd1134 : o_data <= 16'hEB2D;
            12'd1135 : o_data <= 16'hF3CF;
            12'd1136 : o_data <= 16'hF4D3;
            12'd1137 : o_data <= 16'hFD96;
            12'd1138 : o_data <= 16'hEDF6;
            12'd1139 : o_data <= 16'hD697;
            12'd1140 : o_data <= 16'hCEB8;
            12'd1141 : o_data <= 16'hDEB9;
            12'd1142 : o_data <= 16'hE73B;
            12'd1143 : o_data <= 16'hD698;
            12'd1144 : o_data <= 16'hFFFD;
            12'd1145 : o_data <= 16'h62C9;
            12'd1146 : o_data <= 16'h0000;
            12'd1147 : o_data <= 16'h0000;
            12'd1148 : o_data <= 16'h0000;
            12'd1149 : o_data <= 16'h0000;
            12'd1150 : o_data <= 16'h0000;
            12'd1151 : o_data <= 16'h0000;
            12'd1152 : o_data <= 16'h0000;
            12'd1153 : o_data <= 16'h0000;
            12'd1154 : o_data <= 16'h0000;
            12'd1155 : o_data <= 16'h0000;
            12'd1156 : o_data <= 16'h0000;
            12'd1157 : o_data <= 16'h0000;
            12'd1158 : o_data <= 16'h2945;
            12'd1159 : o_data <= 16'hFD55;
            12'd1160 : o_data <= 16'hFC71;
            12'd1161 : o_data <= 16'hF3CF;
            12'd1162 : o_data <= 16'hEAEC;
            12'd1163 : o_data <= 16'hF410;
            12'd1164 : o_data <= 16'hF411;
            12'd1165 : o_data <= 16'hF36E;
            12'd1166 : o_data <= 16'hEB2D;
            12'd1167 : o_data <= 16'hF32D;
            12'd1168 : o_data <= 16'hEACC;
            12'd1169 : o_data <= 16'hF2EC;
            12'd1170 : o_data <= 16'hF34E;
            12'd1171 : o_data <= 16'hF36E;
            12'd1172 : o_data <= 16'hEB0D;
            12'd1173 : o_data <= 16'hF30C;
            12'd1174 : o_data <= 16'hF32E;
            12'd1175 : o_data <= 16'hEB2D;
            12'd1176 : o_data <= 16'hF3AF;
            12'd1177 : o_data <= 16'hEA8B;
            12'd1178 : o_data <= 16'hEA8A;
            12'd1179 : o_data <= 16'hF2AC;
            12'd1180 : o_data <= 16'hEB0C;
            12'd1181 : o_data <= 16'hF30D;
            12'd1182 : o_data <= 16'hEB2D;
            12'd1183 : o_data <= 16'hF34D;
            12'd1184 : o_data <= 16'hEB6E;
            12'd1185 : o_data <= 16'hF3CF;
            12'd1186 : o_data <= 16'hF4D3;
            12'd1187 : o_data <= 16'hFD76;
            12'd1188 : o_data <= 16'hEDF6;
            12'd1189 : o_data <= 16'hC656;
            12'd1190 : o_data <= 16'hD6B8;
            12'd1191 : o_data <= 16'hF77B;
            12'd1192 : o_data <= 16'h632B;
            12'd1193 : o_data <= 16'h0000;
            12'd1194 : o_data <= 16'h0000;
            12'd1195 : o_data <= 16'h0000;
            12'd1196 : o_data <= 16'h0000;
            12'd1197 : o_data <= 16'h0000;
            12'd1198 : o_data <= 16'h0000;
            12'd1199 : o_data <= 16'h0000;
            12'd1200 : o_data <= 16'h0000;
            12'd1201 : o_data <= 16'h0000;
            12'd1202 : o_data <= 16'h0000;
            12'd1203 : o_data <= 16'h0000;
            12'd1204 : o_data <= 16'h0000;
            12'd1205 : o_data <= 16'h0000;
            12'd1206 : o_data <= 16'hFE18;
            12'd1207 : o_data <= 16'hFB6E;
            12'd1208 : o_data <= 16'hF2EC;
            12'd1209 : o_data <= 16'hF2AB;
            12'd1210 : o_data <= 16'hF493;
            12'd1211 : o_data <= 16'hF30C;
            12'd1212 : o_data <= 16'hEAEC;
            12'd1213 : o_data <= 16'hEB4E;
            12'd1214 : o_data <= 16'hEB4E;
            12'd1215 : o_data <= 16'hEC32;
            12'd1216 : o_data <= 16'hF4F4;
            12'd1217 : o_data <= 16'hEBAF;
            12'd1218 : o_data <= 16'hEA8B;
            12'd1219 : o_data <= 16'hF24A;
            12'd1220 : o_data <= 16'hEA4A;
            12'd1221 : o_data <= 16'hEA4A;
            12'd1222 : o_data <= 16'hEA4A;
            12'd1223 : o_data <= 16'hF24A;
            12'd1224 : o_data <= 16'hEA6A;
            12'd1225 : o_data <= 16'hF26B;
            12'd1226 : o_data <= 16'hEA6A;
            12'd1227 : o_data <= 16'hEA6A;
            12'd1228 : o_data <= 16'hEA4A;
            12'd1229 : o_data <= 16'hEAAB;
            12'd1230 : o_data <= 16'hF38F;
            12'd1231 : o_data <= 16'hEBCF;
            12'd1232 : o_data <= 16'hF431;
            12'd1233 : o_data <= 16'hF431;
            12'd1234 : o_data <= 16'hF431;
            12'd1235 : o_data <= 16'hF472;
            12'd1236 : o_data <= 16'hF534;
            12'd1237 : o_data <= 16'hFE39;
            12'd1238 : o_data <= 16'h83CD;
            12'd1239 : o_data <= 16'h0000;
            12'd1240 : o_data <= 16'h0000;
            12'd1241 : o_data <= 16'h0000;
            12'd1242 : o_data <= 16'h0000;
            12'd1243 : o_data <= 16'h0000;
            12'd1244 : o_data <= 16'h0000;
            12'd1245 : o_data <= 16'h0000;
            12'd1246 : o_data <= 16'h0000;
            12'd1247 : o_data <= 16'h0000;
            12'd1248 : o_data <= 16'h0000;
            12'd1249 : o_data <= 16'h0000;
            12'd1250 : o_data <= 16'h0000;
            12'd1251 : o_data <= 16'h0000;
            12'd1252 : o_data <= 16'h0000;
            12'd1253 : o_data <= 16'hA451;
            12'd1254 : o_data <= 16'hFACB;
            12'd1255 : o_data <= 16'hF2EC;
            12'd1256 : o_data <= 16'hF28B;
            12'd1257 : o_data <= 16'hF472;
            12'd1258 : o_data <= 16'hF28B;
            12'd1259 : o_data <= 16'hF30D;
            12'd1260 : o_data <= 16'hF30D;
            12'd1261 : o_data <= 16'hF2ED;
            12'd1262 : o_data <= 16'hF515;
            12'd1263 : o_data <= 16'hF493;
            12'd1264 : o_data <= 16'hEBB0;
            12'd1265 : o_data <= 16'hF36F;
            12'd1266 : o_data <= 16'hF32E;
            12'd1267 : o_data <= 16'hEACC;
            12'd1268 : o_data <= 16'hEA4A;
            12'd1269 : o_data <= 16'hF22A;
            12'd1270 : o_data <= 16'hEA29;
            12'd1271 : o_data <= 16'hEA2A;
            12'd1272 : o_data <= 16'hEA09;
            12'd1273 : o_data <= 16'hEA29;
            12'd1274 : o_data <= 16'hF2CC;
            12'd1275 : o_data <= 16'hF411;
            12'd1276 : o_data <= 16'hF3F0;
            12'd1277 : o_data <= 16'hF34E;
            12'd1278 : o_data <= 16'hEA8B;
            12'd1279 : o_data <= 16'hF28B;
            12'd1280 : o_data <= 16'hEAEC;
            12'd1281 : o_data <= 16'hEB2D;
            12'd1282 : o_data <= 16'hF3AE;
            12'd1283 : o_data <= 16'hEBF0;
            12'd1284 : o_data <= 16'hF410;
            12'd1285 : o_data <= 16'hF492;
            12'd1286 : o_data <= 16'hFDF8;
            12'd1287 : o_data <= 16'hE5F6;
            12'd1288 : o_data <= 16'h0000;
            12'd1289 : o_data <= 16'h0000;
            12'd1290 : o_data <= 16'h0000;
            12'd1291 : o_data <= 16'h0000;
            12'd1292 : o_data <= 16'h0000;
            12'd1293 : o_data <= 16'h0000;
            12'd1294 : o_data <= 16'h0000;
            12'd1295 : o_data <= 16'h0000;
            12'd1296 : o_data <= 16'h0000;
            12'd1297 : o_data <= 16'h0000;
            12'd1298 : o_data <= 16'h0000;
            12'd1299 : o_data <= 16'h0000;
            12'd1300 : o_data <= 16'h0000;
            12'd1301 : o_data <= 16'hFD96;
            12'd1302 : o_data <= 16'hFAAB;
            12'd1303 : o_data <= 16'hF34D;
            12'd1304 : o_data <= 16'hFC31;
            12'd1305 : o_data <= 16'hFA8A;
            12'd1306 : o_data <= 16'hF1E9;
            12'd1307 : o_data <= 16'hF26A;
            12'd1308 : o_data <= 16'hF4B3;
            12'd1309 : o_data <= 16'hF492;
            12'd1310 : o_data <= 16'hE9E8;
            12'd1311 : o_data <= 16'hE9E8;
            12'd1312 : o_data <= 16'hEA08;
            12'd1313 : o_data <= 16'hEA08;
            12'd1314 : o_data <= 16'hF1C8;
            12'd1315 : o_data <= 16'hE9E8;
            12'd1316 : o_data <= 16'hF2AB;
            12'd1317 : o_data <= 16'hF2EC;
            12'd1318 : o_data <= 16'hF2ED;
            12'd1319 : o_data <= 16'hF32E;
            12'd1320 : o_data <= 16'hF34E;
            12'd1321 : o_data <= 16'hF32E;
            12'd1322 : o_data <= 16'hEAEC;
            12'd1323 : o_data <= 16'hEA09;
            12'd1324 : o_data <= 16'hEA4A;
            12'd1325 : o_data <= 16'hF2AB;
            12'd1326 : o_data <= 16'hEAAB;
            12'd1327 : o_data <= 16'hEA8B;
            12'd1328 : o_data <= 16'hF28B;
            12'd1329 : o_data <= 16'hEACC;
            12'd1330 : o_data <= 16'hEB0D;
            12'd1331 : o_data <= 16'hF36E;
            12'd1332 : o_data <= 16'hF3EF;
            12'd1333 : o_data <= 16'hF430;
            12'd1334 : o_data <= 16'hF471;
            12'd1335 : o_data <= 16'hFD34;
            12'd1336 : o_data <= 16'hFE59;
            12'd1337 : o_data <= 16'h1082;
            12'd1338 : o_data <= 16'h0000;
            12'd1339 : o_data <= 16'h0000;
            12'd1340 : o_data <= 16'h0000;
            12'd1341 : o_data <= 16'h0000;
            12'd1342 : o_data <= 16'h0000;
            12'd1343 : o_data <= 16'h0000;
            12'd1344 : o_data <= 16'h0000;
            12'd1345 : o_data <= 16'h0000;
            12'd1346 : o_data <= 16'h0000;
            12'd1347 : o_data <= 16'h0000;
            12'd1348 : o_data <= 16'h3186;
            12'd1349 : o_data <= 16'hFBCF;
            12'd1350 : o_data <= 16'hFC73;
            12'd1351 : o_data <= 16'hF36E;
            12'd1352 : o_data <= 16'hE166;
            12'd1353 : o_data <= 16'hD1E8;
            12'd1354 : o_data <= 16'hD36E;
            12'd1355 : o_data <= 16'hCB2C;
            12'd1356 : o_data <= 16'hC945;
            12'd1357 : o_data <= 16'hC125;
            12'd1358 : o_data <= 16'hC186;
            12'd1359 : o_data <= 16'hC166;
            12'd1360 : o_data <= 16'hC966;
            12'd1361 : o_data <= 16'hC104;
            12'd1362 : o_data <= 16'hCA6A;
            12'd1363 : o_data <= 16'hD229;
            12'd1364 : o_data <= 16'hD125;
            12'd1365 : o_data <= 16'hD905;
            12'd1366 : o_data <= 16'hE145;
            12'd1367 : o_data <= 16'hE9A7;
            12'd1368 : o_data <= 16'hF1C8;
            12'd1369 : o_data <= 16'hF208;
            12'd1370 : o_data <= 16'hF209;
            12'd1371 : o_data <= 16'hEA0A;
            12'd1372 : o_data <= 16'hEA4A;
            12'd1373 : o_data <= 16'hEAAC;
            12'd1374 : o_data <= 16'hF32E;
            12'd1375 : o_data <= 16'hF30D;
            12'd1376 : o_data <= 16'hEACC;
            12'd1377 : o_data <= 16'hF2AB;
            12'd1378 : o_data <= 16'hF2AB;
            12'd1379 : o_data <= 16'hEAAB;
            12'd1380 : o_data <= 16'hF34E;
            12'd1381 : o_data <= 16'hEC11;
            12'd1382 : o_data <= 16'hF492;
            12'd1383 : o_data <= 16'hF4F4;
            12'd1384 : o_data <= 16'hFD54;
            12'd1385 : o_data <= 16'hFEBB;
            12'd1386 : o_data <= 16'h10A2;
            12'd1387 : o_data <= 16'h0000;
            12'd1388 : o_data <= 16'h0000;
            12'd1389 : o_data <= 16'h0000;
            12'd1390 : o_data <= 16'h0000;
            12'd1391 : o_data <= 16'h0000;
            12'd1392 : o_data <= 16'h0000;
            12'd1393 : o_data <= 16'h0000;
            12'd1394 : o_data <= 16'h0000;
            12'd1395 : o_data <= 16'h0000;
            12'd1396 : o_data <= 16'h728A;
            12'd1397 : o_data <= 16'hFB8E;
            12'd1398 : o_data <= 16'hD0C3;
            12'd1399 : o_data <= 16'hC125;
            12'd1400 : o_data <= 16'hB905;
            12'd1401 : o_data <= 16'hC1C7;
            12'd1402 : o_data <= 16'hB842;
            12'd1403 : o_data <= 16'hB822;
            12'd1404 : o_data <= 16'hB042;
            12'd1405 : o_data <= 16'hB082;
            12'd1406 : o_data <= 16'hB041;
            12'd1407 : o_data <= 16'hB882;
            12'd1408 : o_data <= 16'hB862;
            12'd1409 : o_data <= 16'hD2EB;
            12'd1410 : o_data <= 16'hB8A2;
            12'd1411 : o_data <= 16'hC0C3;
            12'd1412 : o_data <= 16'hB0E4;
            12'd1413 : o_data <= 16'hC124;
            12'd1414 : o_data <= 16'hB925;
            12'd1415 : o_data <= 16'hC145;
            12'd1416 : o_data <= 16'hC945;
            12'd1417 : o_data <= 16'hD125;
            12'd1418 : o_data <= 16'hD905;
            12'd1419 : o_data <= 16'hF249;
            12'd1420 : o_data <= 16'hFBD0;
            12'd1421 : o_data <= 16'hFBD0;
            12'd1422 : o_data <= 16'hFCB3;
            12'd1423 : o_data <= 16'hF515;
            12'd1424 : o_data <= 16'hFCB3;
            12'd1425 : o_data <= 16'hF431;
            12'd1426 : o_data <= 16'hF3F0;
            12'd1427 : o_data <= 16'hF3AF;
            12'd1428 : o_data <= 16'hF32D;
            12'd1429 : o_data <= 16'hF2CC;
            12'd1430 : o_data <= 16'hF34D;
            12'd1431 : o_data <= 16'hF3CF;
            12'd1432 : o_data <= 16'hF472;
            12'd1433 : o_data <= 16'hFCD2;
            12'd1434 : o_data <= 16'hFDF8;
            12'd1435 : o_data <= 16'h0000;
            12'd1436 : o_data <= 16'h0000;
            12'd1437 : o_data <= 16'h0000;
            12'd1438 : o_data <= 16'h0000;
            12'd1439 : o_data <= 16'h0000;
            12'd1440 : o_data <= 16'h0000;
            12'd1441 : o_data <= 16'h0000;
            12'd1442 : o_data <= 16'h0000;
            12'd1443 : o_data <= 16'h0000;
            12'd1444 : o_data <= 16'h6B0B;
            12'd1445 : o_data <= 16'hF946;
            12'd1446 : o_data <= 16'hC8A4;
            12'd1447 : o_data <= 16'hB082;
            12'd1448 : o_data <= 16'hA186;
            12'd1449 : o_data <= 16'hAB6C;
            12'd1450 : o_data <= 16'h9CB0;
            12'd1451 : o_data <= 16'hADF5;
            12'd1452 : o_data <= 16'hB676;
            12'd1453 : o_data <= 16'hAE15;
            12'd1454 : o_data <= 16'hCEFA;
            12'd1455 : o_data <= 16'hB615;
            12'd1456 : o_data <= 16'hBDB5;
            12'd1457 : o_data <= 16'hB532;
            12'd1458 : o_data <= 16'hB450;
            12'd1459 : o_data <= 16'hAB0A;
            12'd1460 : o_data <= 16'hAA69;
            12'd1461 : o_data <= 16'hA145;
            12'd1462 : o_data <= 16'hA062;
            12'd1463 : o_data <= 16'hB082;
            12'd1464 : o_data <= 16'hC0C3;
            12'd1465 : o_data <= 16'hC104;
            12'd1466 : o_data <= 16'hCA8A;
            12'd1467 : o_data <= 16'hC186;
            12'd1468 : o_data <= 16'hC904;
            12'd1469 : o_data <= 16'hD125;
            12'd1470 : o_data <= 16'hD986;
            12'd1471 : o_data <= 16'hEA8B;
            12'd1472 : o_data <= 16'hF38F;
            12'd1473 : o_data <= 16'hFC32;
            12'd1474 : o_data <= 16'hF3D0;
            12'd1475 : o_data <= 16'hF34E;
            12'd1476 : o_data <= 16'hF30C;
            12'd1477 : o_data <= 16'hF2CC;
            12'd1478 : o_data <= 16'hF2EC;
            12'd1479 : o_data <= 16'hF32D;
            12'd1480 : o_data <= 16'hF3CF;
            12'd1481 : o_data <= 16'hFC92;
            12'd1482 : o_data <= 16'hFCF3;
            12'd1483 : o_data <= 16'h5208;
            12'd1484 : o_data <= 16'h0000;
            12'd1485 : o_data <= 16'h0000;
            12'd1486 : o_data <= 16'h0000;
            12'd1487 : o_data <= 16'h0000;
            12'd1488 : o_data <= 16'h0000;
            12'd1489 : o_data <= 16'h0000;
            12'd1490 : o_data <= 16'h0000;
            12'd1491 : o_data <= 16'h0000;
            12'd1492 : o_data <= 16'h0000;
            12'd1493 : o_data <= 16'hA470;
            12'd1494 : o_data <= 16'hBDB4;
            12'd1495 : o_data <= 16'hD79C;
            12'd1496 : o_data <= 16'hDF9C;
            12'd1497 : o_data <= 16'hEF9D;
            12'd1498 : o_data <= 16'hEF7D;
            12'd1499 : o_data <= 16'hF7BD;
            12'd1500 : o_data <= 16'hEF5D;
            12'd1501 : o_data <= 16'hEF7C;
            12'd1502 : o_data <= 16'hEF7D;
            12'd1503 : o_data <= 16'hEF7D;
            12'd1504 : o_data <= 16'hE73B;
            12'd1505 : o_data <= 16'hE75C;
            12'd1506 : o_data <= 16'hDEFA;
            12'd1507 : o_data <= 16'hE79D;
            12'd1508 : o_data <= 16'hDF9C;
            12'd1509 : o_data <= 16'hDFBD;
            12'd1510 : o_data <= 16'hC719;
            12'd1511 : o_data <= 16'hADD5;
            12'd1512 : o_data <= 16'h9C0E;
            12'd1513 : o_data <= 16'hA2CA;
            12'd1514 : o_data <= 16'hA0A2;
            12'd1515 : o_data <= 16'hB862;
            12'd1516 : o_data <= 16'hC104;
            12'd1517 : o_data <= 16'hC125;
            12'd1518 : o_data <= 16'hC945;
            12'd1519 : o_data <= 16'hC966;
            12'd1520 : o_data <= 16'hD166;
            12'd1521 : o_data <= 16'hE229;
            12'd1522 : o_data <= 16'hFB4E;
            12'd1523 : o_data <= 16'hFBF1;
            12'd1524 : o_data <= 16'hFBD0;
            12'd1525 : o_data <= 16'hF34D;
            12'd1526 : o_data <= 16'hF2EC;
            12'd1527 : o_data <= 16'hFAEC;
            12'd1528 : o_data <= 16'hF32D;
            12'd1529 : o_data <= 16'hF3CF;
            12'd1530 : o_data <= 16'hFC71;
            12'd1531 : o_data <= 16'h9B8E;
            12'd1532 : o_data <= 16'h0000;
            12'd1533 : o_data <= 16'h0000;
            12'd1534 : o_data <= 16'h0000;
            12'd1535 : o_data <= 16'h0000;
            12'd1536 : o_data <= 16'h0000;
            12'd1537 : o_data <= 16'h0000;
            12'd1538 : o_data <= 16'h0000;
            12'd1539 : o_data <= 16'h0000;
            12'd1540 : o_data <= 16'h0000;
            12'd1541 : o_data <= 16'h634C;
            12'd1542 : o_data <= 16'hEF7C;
            12'd1543 : o_data <= 16'hF7BE;
            12'd1544 : o_data <= 16'hEF9D;
            12'd1545 : o_data <= 16'hF79D;
            12'd1546 : o_data <= 16'hE75C;
            12'd1547 : o_data <= 16'hDEFA;
            12'd1548 : o_data <= 16'hE73B;
            12'd1549 : o_data <= 16'hE71B;
            12'd1550 : o_data <= 16'hEF5C;
            12'd1551 : o_data <= 16'hE73B;
            12'd1552 : o_data <= 16'hE71B;
            12'd1553 : o_data <= 16'hEF9D;
            12'd1554 : o_data <= 16'hF79D;
            12'd1555 : o_data <= 16'hEF7D;
            12'd1556 : o_data <= 16'hEF7D;
            12'd1557 : o_data <= 16'hE6FA;
            12'd1558 : o_data <= 16'hEF9D;
            12'd1559 : o_data <= 16'hEF5B;
            12'd1560 : o_data <= 16'hE75C;
            12'd1561 : o_data <= 16'hDF3B;
            12'd1562 : o_data <= 16'hE7FE;
            12'd1563 : o_data <= 16'hAD94;
            12'd1564 : o_data <= 16'hA32B;
            12'd1565 : o_data <= 16'h9861;
            12'd1566 : o_data <= 16'hC0A3;
            12'd1567 : o_data <= 16'hC104;
            12'd1568 : o_data <= 16'hC965;
            12'd1569 : o_data <= 16'hD167;
            12'd1570 : o_data <= 16'hD145;
            12'd1571 : o_data <= 16'hE1A7;
            12'd1572 : o_data <= 16'hFAEC;
            12'd1573 : o_data <= 16'hFB8F;
            12'd1574 : o_data <= 16'hFB0D;
            12'd1575 : o_data <= 16'hF2CC;
            12'd1576 : o_data <= 16'hFAEC;
            12'd1577 : o_data <= 16'hF34D;
            12'd1578 : o_data <= 16'hFC51;
            12'd1579 : o_data <= 16'h9BCF;
            12'd1580 : o_data <= 16'h0000;
            12'd1581 : o_data <= 16'h0000;
            12'd1582 : o_data <= 16'h0000;
            12'd1583 : o_data <= 16'h0000;
            12'd1584 : o_data <= 16'h0000;
            12'd1585 : o_data <= 16'h0000;
            12'd1586 : o_data <= 16'h0000;
            12'd1587 : o_data <= 16'h0000;
            12'd1588 : o_data <= 16'h0000;
            12'd1589 : o_data <= 16'h10A2;
            12'd1590 : o_data <= 16'hFFFF;
            12'd1591 : o_data <= 16'hDEFA;
            12'd1592 : o_data <= 16'hDEFA;
            12'd1593 : o_data <= 16'hEF5C;
            12'd1594 : o_data <= 16'hE75B;
            12'd1595 : o_data <= 16'hE73B;
            12'd1596 : o_data <= 16'hE73B;
            12'd1597 : o_data <= 16'hDEFA;
            12'd1598 : o_data <= 16'hD6B9;
            12'd1599 : o_data <= 16'hD6D9;
            12'd1600 : o_data <= 16'hEF5C;
            12'd1601 : o_data <= 16'hE71A;
            12'd1602 : o_data <= 16'hDF1B;
            12'd1603 : o_data <= 16'hE73B;
            12'd1604 : o_data <= 16'hE73B;
            12'd1605 : o_data <= 16'hE73B;
            12'd1606 : o_data <= 16'hE73C;
            12'd1607 : o_data <= 16'hEF5C;
            12'd1608 : o_data <= 16'hEF7D;
            12'd1609 : o_data <= 16'hEF7D;
            12'd1610 : o_data <= 16'hEF7D;
            12'd1611 : o_data <= 16'hEF9C;
            12'd1612 : o_data <= 16'hEFBD;
            12'd1613 : o_data <= 16'hDFBD;
            12'd1614 : o_data <= 16'hA4F2;
            12'd1615 : o_data <= 16'hA185;
            12'd1616 : o_data <= 16'hB862;
            12'd1617 : o_data <= 16'hC0E3;
            12'd1618 : o_data <= 16'hCA29;
            12'd1619 : o_data <= 16'hD2AB;
            12'd1620 : o_data <= 16'hD1A7;
            12'd1621 : o_data <= 16'hEA29;
            12'd1622 : o_data <= 16'hFB4D;
            12'd1623 : o_data <= 16'hFBAF;
            12'd1624 : o_data <= 16'hFBAF;
            12'd1625 : o_data <= 16'hFC72;
            12'd1626 : o_data <= 16'hFB8E;
            12'd1627 : o_data <= 16'h7B6D;
            12'd1628 : o_data <= 16'h0000;
            12'd1629 : o_data <= 16'h0000;
            12'd1630 : o_data <= 16'h0000;
            12'd1631 : o_data <= 16'h0000;
            12'd1632 : o_data <= 16'h0000;
            12'd1633 : o_data <= 16'h0000;
            12'd1634 : o_data <= 16'h0000;
            12'd1635 : o_data <= 16'h0000;
            12'd1636 : o_data <= 16'h0000;
            12'd1637 : o_data <= 16'h0000;
            12'd1638 : o_data <= 16'h630A;
            12'd1639 : o_data <= 16'hE719;
            12'd1640 : o_data <= 16'hD6D9;
            12'd1641 : o_data <= 16'hDEDA;
            12'd1642 : o_data <= 16'hC657;
            12'd1643 : o_data <= 16'hD698;
            12'd1644 : o_data <= 16'hD6B9;
            12'd1645 : o_data <= 16'hD698;
            12'd1646 : o_data <= 16'hD6B9;
            12'd1647 : o_data <= 16'hE71B;
            12'd1648 : o_data <= 16'hCE77;
            12'd1649 : o_data <= 16'hDEFA;
            12'd1650 : o_data <= 16'hDEDA;
            12'd1651 : o_data <= 16'hD6B9;
            12'd1652 : o_data <= 16'hE71B;
            12'd1653 : o_data <= 16'hDF1B;
            12'd1654 : o_data <= 16'hDEFA;
            12'd1655 : o_data <= 16'hDF1A;
            12'd1656 : o_data <= 16'hE73C;
            12'd1657 : o_data <= 16'hEF7C;
            12'd1658 : o_data <= 16'hEF7C;
            12'd1659 : o_data <= 16'hF7BE;
            12'd1660 : o_data <= 16'hEF7D;
            12'd1661 : o_data <= 16'hEF9D;
            12'd1662 : o_data <= 16'hE75B;
            12'd1663 : o_data <= 16'hD75B;
            12'd1664 : o_data <= 16'hA5B4;
            12'd1665 : o_data <= 16'h91A6;
            12'd1666 : o_data <= 16'hC125;
            12'd1667 : o_data <= 16'hC0C3;
            12'd1668 : o_data <= 16'hC925;
            12'd1669 : o_data <= 16'hC8E5;
            12'd1670 : o_data <= 16'hE105;
            12'd1671 : o_data <= 16'hFA29;
            12'd1672 : o_data <= 16'hFB4D;
            12'd1673 : o_data <= 16'hFB8E;
            12'd1674 : o_data <= 16'hFB6E;
            12'd1675 : o_data <= 16'h4249;
            12'd1676 : o_data <= 16'h0000;
            12'd1677 : o_data <= 16'h0000;
            12'd1678 : o_data <= 16'h0000;
            12'd1679 : o_data <= 16'h0000;
            12'd1680 : o_data <= 16'h0000;
            12'd1681 : o_data <= 16'h0000;
            12'd1682 : o_data <= 16'h0000;
            12'd1683 : o_data <= 16'h0000;
            12'd1684 : o_data <= 16'h0000;
            12'd1685 : o_data <= 16'h0000;
            12'd1686 : o_data <= 16'h0000;
            12'd1687 : o_data <= 16'h39C6;
            12'd1688 : o_data <= 16'hBE15;
            12'd1689 : o_data <= 16'hD677;
            12'd1690 : o_data <= 16'hE73B;
            12'd1691 : o_data <= 16'hDEFA;
            12'd1692 : o_data <= 16'hDEDA;
            12'd1693 : o_data <= 16'hD6D9;
            12'd1694 : o_data <= 16'hD6D9;
            12'd1695 : o_data <= 16'hCE78;
            12'd1696 : o_data <= 16'hC657;
            12'd1697 : o_data <= 16'hDEFA;
            12'd1698 : o_data <= 16'hCE78;
            12'd1699 : o_data <= 16'hCE77;
            12'd1700 : o_data <= 16'hE71B;
            12'd1701 : o_data <= 16'hCE98;
            12'd1702 : o_data <= 16'hE71B;
            12'd1703 : o_data <= 16'hDEFA;
            12'd1704 : o_data <= 16'hDF1A;
            12'd1705 : o_data <= 16'hDEFA;
            12'd1706 : o_data <= 16'hEF5C;
            12'd1707 : o_data <= 16'hE71B;
            12'd1708 : o_data <= 16'hE73B;
            12'd1709 : o_data <= 16'hE73C;
            12'd1710 : o_data <= 16'hE71B;
            12'd1711 : o_data <= 16'hF7BE;
            12'd1712 : o_data <= 16'hEF7D;
            12'd1713 : o_data <= 16'hE7DD;
            12'd1714 : o_data <= 16'hA552;
            12'd1715 : o_data <= 16'hA145;
            12'd1716 : o_data <= 16'hB882;
            12'd1717 : o_data <= 16'hC145;
            12'd1718 : o_data <= 16'hC105;
            12'd1719 : o_data <= 16'hD105;
            12'd1720 : o_data <= 16'hE905;
            12'd1721 : o_data <= 16'hF966;
            12'd1722 : o_data <= 16'hFD35;
            12'd1723 : o_data <= 16'h0000;
            12'd1724 : o_data <= 16'h0000;
            12'd1725 : o_data <= 16'h0000;
            12'd1726 : o_data <= 16'h0000;
            12'd1727 : o_data <= 16'h0000;
            12'd1728 : o_data <= 16'h0000;
            12'd1729 : o_data <= 16'h0000;
            12'd1730 : o_data <= 16'h0000;
            12'd1731 : o_data <= 16'h0000;
            12'd1732 : o_data <= 16'h0000;
            12'd1733 : o_data <= 16'h0000;
            12'd1734 : o_data <= 16'h0000;
            12'd1735 : o_data <= 16'h0000;
            12'd1736 : o_data <= 16'h0000;
            12'd1737 : o_data <= 16'h18C2;
            12'd1738 : o_data <= 16'h632B;
            12'd1739 : o_data <= 16'hAD93;
            12'd1740 : o_data <= 16'hF79C;
            12'd1741 : o_data <= 16'hDED9;
            12'd1742 : o_data <= 16'hCE57;
            12'd1743 : o_data <= 16'hDED9;
            12'd1744 : o_data <= 16'hD6B9;
            12'd1745 : o_data <= 16'hCE57;
            12'd1746 : o_data <= 16'hCE78;
            12'd1747 : o_data <= 16'hDEFA;
            12'd1748 : o_data <= 16'hDED9;
            12'd1749 : o_data <= 16'hBDF5;
            12'd1750 : o_data <= 16'hE71B;
            12'd1751 : o_data <= 16'hDEFA;
            12'd1752 : o_data <= 16'hD698;
            12'd1753 : o_data <= 16'hE71A;
            12'd1754 : o_data <= 16'hDF1A;
            12'd1755 : o_data <= 16'hCE98;
            12'd1756 : o_data <= 16'hDF1B;
            12'd1757 : o_data <= 16'hDED9;
            12'd1758 : o_data <= 16'hE73B;
            12'd1759 : o_data <= 16'hE75C;
            12'd1760 : o_data <= 16'hF79D;
            12'd1761 : o_data <= 16'hE73B;
            12'd1762 : o_data <= 16'hF7BE;
            12'd1763 : o_data <= 16'hDFDD;
            12'd1764 : o_data <= 16'hACD1;
            12'd1765 : o_data <= 16'hA0C3;
            12'd1766 : o_data <= 16'hA8A3;
            12'd1767 : o_data <= 16'hA8E3;
            12'd1768 : o_data <= 16'hB0E4;
            12'd1769 : o_data <= 16'hE0C4;
            12'd1770 : o_data <= 16'hA451;
            12'd1771 : o_data <= 16'h0000;
            12'd1772 : o_data <= 16'h0000;
            12'd1773 : o_data <= 16'h0000;
            12'd1774 : o_data <= 16'h0000;
            12'd1775 : o_data <= 16'h0000;
            12'd1776 : o_data <= 16'h0000;
            12'd1777 : o_data <= 16'h0000;
            12'd1778 : o_data <= 16'h0000;
            12'd1779 : o_data <= 16'h0000;
            12'd1780 : o_data <= 16'h0000;
            12'd1781 : o_data <= 16'h0000;
            12'd1782 : o_data <= 16'h0000;
            12'd1783 : o_data <= 16'h0000;
            12'd1784 : o_data <= 16'h0000;
            12'd1785 : o_data <= 16'h0000;
            12'd1786 : o_data <= 16'h0000;
            12'd1787 : o_data <= 16'h0000;
            12'd1788 : o_data <= 16'h0000;
            12'd1789 : o_data <= 16'h3A07;
            12'd1790 : o_data <= 16'h7BEE;
            12'd1791 : o_data <= 16'hC616;
            12'd1792 : o_data <= 16'hDEF9;
            12'd1793 : o_data <= 16'hCE77;
            12'd1794 : o_data <= 16'hD6B8;
            12'd1795 : o_data <= 16'hCE98;
            12'd1796 : o_data <= 16'hDEB9;
            12'd1797 : o_data <= 16'hE73B;
            12'd1798 : o_data <= 16'hDED9;
            12'd1799 : o_data <= 16'hCE98;
            12'd1800 : o_data <= 16'hEF3C;
            12'd1801 : o_data <= 16'hCE98;
            12'd1802 : o_data <= 16'hD6B9;
            12'd1803 : o_data <= 16'hD6B9;
            12'd1804 : o_data <= 16'hDED9;
            12'd1805 : o_data <= 16'hDEDA;
            12'd1806 : o_data <= 16'hCE77;
            12'd1807 : o_data <= 16'hDEFB;
            12'd1808 : o_data <= 16'hDEFA;
            12'd1809 : o_data <= 16'hDF1A;
            12'd1810 : o_data <= 16'hEF5C;
            12'd1811 : o_data <= 16'hE71B;
            12'd1812 : o_data <= 16'hEF9D;
            12'd1813 : o_data <= 16'hD79C;
            12'd1814 : o_data <= 16'hACB0;
            12'd1815 : o_data <= 16'h9A28;
            12'd1816 : o_data <= 16'hBA8A;
            12'd1817 : o_data <= 16'hDD13;
            12'd1818 : o_data <= 16'h0000;
            12'd1819 : o_data <= 16'h0000;
            12'd1820 : o_data <= 16'h0000;
            12'd1821 : o_data <= 16'h0000;
            12'd1822 : o_data <= 16'h0000;
            12'd1823 : o_data <= 16'h0000;
            12'd1824 : o_data <= 16'h0000;
            12'd1825 : o_data <= 16'h0000;
            12'd1826 : o_data <= 16'h0000;
            12'd1827 : o_data <= 16'h0000;
            12'd1828 : o_data <= 16'h0000;
            12'd1829 : o_data <= 16'h0000;
            12'd1830 : o_data <= 16'h0000;
            12'd1831 : o_data <= 16'h0000;
            12'd1832 : o_data <= 16'h0000;
            12'd1833 : o_data <= 16'h0000;
            12'd1834 : o_data <= 16'h0000;
            12'd1835 : o_data <= 16'h0000;
            12'd1836 : o_data <= 16'h0000;
            12'd1837 : o_data <= 16'h0000;
            12'd1838 : o_data <= 16'h0000;
            12'd1839 : o_data <= 16'h0000;
            12'd1840 : o_data <= 16'h0000;
            12'd1841 : o_data <= 16'h4227;
            12'd1842 : o_data <= 16'h632B;
            12'd1843 : o_data <= 16'h8C4F;
            12'd1844 : o_data <= 16'hC636;
            12'd1845 : o_data <= 16'hDEF9;
            12'd1846 : o_data <= 16'hD698;
            12'd1847 : o_data <= 16'hDEF9;
            12'd1848 : o_data <= 16'hBE16;
            12'd1849 : o_data <= 16'hD6B9;
            12'd1850 : o_data <= 16'hD6B8;
            12'd1851 : o_data <= 16'hC616;
            12'd1852 : o_data <= 16'hBDD5;
            12'd1853 : o_data <= 16'hCE77;
            12'd1854 : o_data <= 16'hDEFA;
            12'd1855 : o_data <= 16'hD698;
            12'd1856 : o_data <= 16'hD6B9;
            12'd1857 : o_data <= 16'hD698;
            12'd1858 : o_data <= 16'hDF1B;
            12'd1859 : o_data <= 16'hE71B;
            12'd1860 : o_data <= 16'hDF1B;
            12'd1861 : o_data <= 16'hEF7C;
            12'd1862 : o_data <= 16'hD6FA;
            12'd1863 : o_data <= 16'hEF9D;
            12'd1864 : o_data <= 16'hADF5;
            12'd1865 : o_data <= 16'h0000;
            12'd1866 : o_data <= 16'h0000;
            12'd1867 : o_data <= 16'h0000;
            12'd1868 : o_data <= 16'h0000;
            12'd1869 : o_data <= 16'h0000;
            12'd1870 : o_data <= 16'h0000;
            12'd1871 : o_data <= 16'h0000;
            12'd1872 : o_data <= 16'h0000;
            12'd1873 : o_data <= 16'h0000;
            12'd1874 : o_data <= 16'h0000;
            12'd1875 : o_data <= 16'h0000;
            12'd1876 : o_data <= 16'h0000;
            12'd1877 : o_data <= 16'h0000;
            12'd1878 : o_data <= 16'h0000;
            12'd1879 : o_data <= 16'h0000;
            12'd1880 : o_data <= 16'h0000;
            12'd1881 : o_data <= 16'h0000;
            12'd1882 : o_data <= 16'h0000;
            12'd1883 : o_data <= 16'h0000;
            12'd1884 : o_data <= 16'h0000;
            12'd1885 : o_data <= 16'h0000;
            12'd1886 : o_data <= 16'h0000;
            12'd1887 : o_data <= 16'h0000;
            12'd1888 : o_data <= 16'h0000;
            12'd1889 : o_data <= 16'h0000;
            12'd1890 : o_data <= 16'h0000;
            12'd1891 : o_data <= 16'h0000;
            12'd1892 : o_data <= 16'h0000;
            12'd1893 : o_data <= 16'h0000;
            12'd1894 : o_data <= 16'h2123;
            12'd1895 : o_data <= 16'h7BCE;
            12'd1896 : o_data <= 16'hDEF9;
            12'd1897 : o_data <= 16'hCE97;
            12'd1898 : o_data <= 16'hDED9;
            12'd1899 : o_data <= 16'hE73A;
            12'd1900 : o_data <= 16'hDF3B;
            12'd1901 : o_data <= 16'hD6B9;
            12'd1902 : o_data <= 16'hCE98;
            12'd1903 : o_data <= 16'hD698;
            12'd1904 : o_data <= 16'hD698;
            12'd1905 : o_data <= 16'hD6B9;
            12'd1906 : o_data <= 16'hC636;
            12'd1907 : o_data <= 16'hE71B;
            12'd1908 : o_data <= 16'hCE77;
            12'd1909 : o_data <= 16'hD6B9;
            12'd1910 : o_data <= 16'hF79D;
            12'd1911 : o_data <= 16'hFFFE;
            12'd1912 : o_data <= 16'h0040;
            12'd1913 : o_data <= 16'h0000;
            12'd1914 : o_data <= 16'h0000;
            12'd1915 : o_data <= 16'h0000;
            12'd1916 : o_data <= 16'h0000;
            12'd1917 : o_data <= 16'h0000;
            12'd1918 : o_data <= 16'h0000;
            12'd1919 : o_data <= 16'h0000;
            12'd1920 : o_data <= 16'h0000;
            12'd1921 : o_data <= 16'h0000;
            12'd1922 : o_data <= 16'h0000;
            12'd1923 : o_data <= 16'h0000;
            12'd1924 : o_data <= 16'h0000;
            12'd1925 : o_data <= 16'h0000;
            12'd1926 : o_data <= 16'h0000;
            12'd1927 : o_data <= 16'h0000;
            12'd1928 : o_data <= 16'h0000;
            12'd1929 : o_data <= 16'h0000;
            12'd1930 : o_data <= 16'h0000;
            12'd1931 : o_data <= 16'h0000;
            12'd1932 : o_data <= 16'h0000;
            12'd1933 : o_data <= 16'h0000;
            12'd1934 : o_data <= 16'h0000;
            12'd1935 : o_data <= 16'h0000;
            12'd1936 : o_data <= 16'h0000;
            12'd1937 : o_data <= 16'h0000;
            12'd1938 : o_data <= 16'h0000;
            12'd1939 : o_data <= 16'h0000;
            12'd1940 : o_data <= 16'h0000;
            12'd1941 : o_data <= 16'h0000;
            12'd1942 : o_data <= 16'h0000;
            12'd1943 : o_data <= 16'h0000;
            12'd1944 : o_data <= 16'h0000;
            12'd1945 : o_data <= 16'h0000;
            12'd1946 : o_data <= 16'h0000;
            12'd1947 : o_data <= 16'h39C6;
            12'd1948 : o_data <= 16'h52A9;
            12'd1949 : o_data <= 16'h5AA9;
            12'd1950 : o_data <= 16'h8C4F;
            12'd1951 : o_data <= 16'hD6B9;
            12'd1952 : o_data <= 16'hD6D8;
            12'd1953 : o_data <= 16'hDED9;
            12'd1954 : o_data <= 16'hD6F9;
            12'd1955 : o_data <= 16'hD6B8;
            12'd1956 : o_data <= 16'hC616;
            12'd1957 : o_data <= 16'hDED9;
            12'd1958 : o_data <= 16'h9D11;
            12'd1959 : o_data <= 16'h0861;
            12'd1960 : o_data <= 16'h0000;
            12'd1961 : o_data <= 16'h0000;
            12'd1962 : o_data <= 16'h0000;
            12'd1963 : o_data <= 16'h0000;
            12'd1964 : o_data <= 16'h0000;
            12'd1965 : o_data <= 16'h0000;
            12'd1966 : o_data <= 16'h0000;
            12'd1967 : o_data <= 16'h0000;
            12'd1968 : o_data <= 16'h0000;
            12'd1969 : o_data <= 16'h0000;
            12'd1970 : o_data <= 16'h0000;
            12'd1971 : o_data <= 16'h0000;
            12'd1972 : o_data <= 16'h0000;
            12'd1973 : o_data <= 16'h0000;
            12'd1974 : o_data <= 16'h0000;
            12'd1975 : o_data <= 16'h0000;
            12'd1976 : o_data <= 16'h0000;
            12'd1977 : o_data <= 16'h0000;
            12'd1978 : o_data <= 16'h0000;
            12'd1979 : o_data <= 16'h0000;
            12'd1980 : o_data <= 16'h0000;
            12'd1981 : o_data <= 16'h0000;
            12'd1982 : o_data <= 16'h0000;
            12'd1983 : o_data <= 16'h0000;
            12'd1984 : o_data <= 16'h0000;
            12'd1985 : o_data <= 16'h0000;
            12'd1986 : o_data <= 16'h0000;
            12'd1987 : o_data <= 16'h0000;
            12'd1988 : o_data <= 16'h0000;
            12'd1989 : o_data <= 16'h0000;
            12'd1990 : o_data <= 16'h0000;
            12'd1991 : o_data <= 16'h0000;
            12'd1992 : o_data <= 16'h0000;
            12'd1993 : o_data <= 16'h0000;
            12'd1994 : o_data <= 16'h0000;
            12'd1995 : o_data <= 16'h0000;
            12'd1996 : o_data <= 16'h0000;
            12'd1997 : o_data <= 16'h0000;
            12'd1998 : o_data <= 16'h0000;
            12'd1999 : o_data <= 16'h0000;
            12'd2000 : o_data <= 16'h0000;
            12'd2001 : o_data <= 16'h0000;
            12'd2002 : o_data <= 16'h0840;
            12'd2003 : o_data <= 16'h4A48;
            12'd2004 : o_data <= 16'h52CA;
            12'd2005 : o_data <= 16'h0000;
            12'd2006 : o_data <= 16'h0000;
            12'd2007 : o_data <= 16'h0000;
            12'd2008 : o_data <= 16'h0000;
            12'd2009 : o_data <= 16'h0000;
            12'd2010 : o_data <= 16'h0000;
            12'd2011 : o_data <= 16'h0000;
            12'd2012 : o_data <= 16'h0000;
            12'd2013 : o_data <= 16'h0000;
            12'd2014 : o_data <= 16'h0000;
            12'd2015 : o_data <= 16'h0000;
            12'd2016 : o_data <= 16'h0000;
            12'd2017 : o_data <= 16'h0000;
            12'd2018 : o_data <= 16'h0000;
            12'd2019 : o_data <= 16'h0000;
            12'd2020 : o_data <= 16'h0000;
            12'd2021 : o_data <= 16'h0000;
            12'd2022 : o_data <= 16'h0000;
            12'd2023 : o_data <= 16'h0000;
            12'd2024 : o_data <= 16'h0000;
            12'd2025 : o_data <= 16'h0000;
            12'd2026 : o_data <= 16'h0000;
            12'd2027 : o_data <= 16'h0000;
            12'd2028 : o_data <= 16'h0000;
            12'd2029 : o_data <= 16'h0000;
            12'd2030 : o_data <= 16'h0000;
            12'd2031 : o_data <= 16'h0000;
            12'd2032 : o_data <= 16'h0000;
            12'd2033 : o_data <= 16'h0000;
            12'd2034 : o_data <= 16'h0000;
            12'd2035 : o_data <= 16'h0000;
            12'd2036 : o_data <= 16'h0000;
            12'd2037 : o_data <= 16'h0000;
            12'd2038 : o_data <= 16'h0000;
            12'd2039 : o_data <= 16'h0000;
            12'd2040 : o_data <= 16'h0000;
            12'd2041 : o_data <= 16'h0000;
            12'd2042 : o_data <= 16'h0000;
            12'd2043 : o_data <= 16'h0000;
            12'd2044 : o_data <= 16'h0000;
            12'd2045 : o_data <= 16'h0000;
            12'd2046 : o_data <= 16'h0000;
            12'd2047 : o_data <= 16'h0000;
            12'd2048 : o_data <= 16'h0000;
            12'd2049 : o_data <= 16'h0000;
            12'd2050 : o_data <= 16'h0000;
            12'd2051 : o_data <= 16'h0000;
            12'd2052 : o_data <= 16'h0000;
            12'd2053 : o_data <= 16'h0000;
            12'd2054 : o_data <= 16'h0000;
            12'd2055 : o_data <= 16'h0000;
            12'd2056 : o_data <= 16'h0000;
            12'd2057 : o_data <= 16'h0000;
            12'd2058 : o_data <= 16'h0000;
            12'd2059 : o_data <= 16'h0000;
            12'd2060 : o_data <= 16'h0000;
            12'd2061 : o_data <= 16'h0000;
            12'd2062 : o_data <= 16'h0000;
            12'd2063 : o_data <= 16'h0000;
            12'd2064 : o_data <= 16'h0000;
            12'd2065 : o_data <= 16'h0000;
            12'd2066 : o_data <= 16'h0000;
            12'd2067 : o_data <= 16'h0000;
            12'd2068 : o_data <= 16'h0000;
            12'd2069 : o_data <= 16'h0000;
            12'd2070 : o_data <= 16'h0000;
            12'd2071 : o_data <= 16'h0000;
            12'd2072 : o_data <= 16'h0000;
            12'd2073 : o_data <= 16'h0000;
            12'd2074 : o_data <= 16'h0000;
            12'd2075 : o_data <= 16'h0000;
            12'd2076 : o_data <= 16'h0000;
            12'd2077 : o_data <= 16'h0000;
            12'd2078 : o_data <= 16'h0000;
            12'd2079 : o_data <= 16'h0000;
            12'd2080 : o_data <= 16'h0000;
            12'd2081 : o_data <= 16'h0000;
            12'd2082 : o_data <= 16'h0000;
            12'd2083 : o_data <= 16'h0000;
            12'd2084 : o_data <= 16'h0000;
            12'd2085 : o_data <= 16'h0000;
            12'd2086 : o_data <= 16'h0000;
            12'd2087 : o_data <= 16'h0000;
            12'd2088 : o_data <= 16'h0000;
            12'd2089 : o_data <= 16'h0000;
            12'd2090 : o_data <= 16'h0000;
            12'd2091 : o_data <= 16'h0000;
            12'd2092 : o_data <= 16'h0000;
            12'd2093 : o_data <= 16'h0000;
            12'd2094 : o_data <= 16'h0000;
            12'd2095 : o_data <= 16'h0000;
            12'd2096 : o_data <= 16'h0000;
            12'd2097 : o_data <= 16'h0000;
            12'd2098 : o_data <= 16'h0000;
            12'd2099 : o_data <= 16'h0000;
            12'd2100 : o_data <= 16'h0000;
            12'd2101 : o_data <= 16'h0000;
            12'd2102 : o_data <= 16'h0000;
            12'd2103 : o_data <= 16'h0000;
            12'd2104 : o_data <= 16'h0000;
            12'd2105 : o_data <= 16'h0000;
            12'd2106 : o_data <= 16'h0000;
            12'd2107 : o_data <= 16'h0000;
            12'd2108 : o_data <= 16'h0000;
            12'd2109 : o_data <= 16'h0000;
            12'd2110 : o_data <= 16'h0000;
            12'd2111 : o_data <= 16'h0000;
            12'd2112 : o_data <= 16'h0000;
            12'd2113 : o_data <= 16'h0000;
            12'd2114 : o_data <= 16'h0000;
            12'd2115 : o_data <= 16'h0000;
            12'd2116 : o_data <= 16'h0000;
            12'd2117 : o_data <= 16'h0000;
            12'd2118 : o_data <= 16'h0000;
            12'd2119 : o_data <= 16'h0000;
            12'd2120 : o_data <= 16'h0000;
            12'd2121 : o_data <= 16'h0000;
            12'd2122 : o_data <= 16'h0000;
            12'd2123 : o_data <= 16'h0000;
            12'd2124 : o_data <= 16'h0000;
            12'd2125 : o_data <= 16'h0000;
            12'd2126 : o_data <= 16'h0000;
            12'd2127 : o_data <= 16'h0000;
            12'd2128 : o_data <= 16'h0000;
            12'd2129 : o_data <= 16'h0000;
            12'd2130 : o_data <= 16'h0000;
            12'd2131 : o_data <= 16'h0000;
            12'd2132 : o_data <= 16'h0000;
            12'd2133 : o_data <= 16'h0000;
            12'd2134 : o_data <= 16'h0000;
            12'd2135 : o_data <= 16'h0000;
            12'd2136 : o_data <= 16'h0000;
            12'd2137 : o_data <= 16'h0000;
            12'd2138 : o_data <= 16'h0000;
            12'd2139 : o_data <= 16'h0000;
            12'd2140 : o_data <= 16'h0000;
            12'd2141 : o_data <= 16'h0000;
            12'd2142 : o_data <= 16'h0000;
            12'd2143 : o_data <= 16'h0000;
            12'd2144 : o_data <= 16'h0000;
            12'd2145 : o_data <= 16'h0000;
            12'd2146 : o_data <= 16'h0000;
            12'd2147 : o_data <= 16'h0000;
            12'd2148 : o_data <= 16'h0000;
            12'd2149 : o_data <= 16'h0000;
            12'd2150 : o_data <= 16'h0000;
            12'd2151 : o_data <= 16'h0000;
            12'd2152 : o_data <= 16'h0000;
            12'd2153 : o_data <= 16'h0000;
            12'd2154 : o_data <= 16'h0000;
            12'd2155 : o_data <= 16'h0000;
            12'd2156 : o_data <= 16'h0000;
            12'd2157 : o_data <= 16'h0000;
            12'd2158 : o_data <= 16'h0000;
            12'd2159 : o_data <= 16'h0000;
            12'd2160 : o_data <= 16'h0000;
            12'd2161 : o_data <= 16'h0000;
            12'd2162 : o_data <= 16'h0000;
            12'd2163 : o_data <= 16'h0000;
            12'd2164 : o_data <= 16'h0000;
            12'd2165 : o_data <= 16'h0000;
            12'd2166 : o_data <= 16'h0000;
            12'd2167 : o_data <= 16'h0000;
            12'd2168 : o_data <= 16'h0000;
            12'd2169 : o_data <= 16'h0000;
            12'd2170 : o_data <= 16'h0000;
            12'd2171 : o_data <= 16'h0000;
            12'd2172 : o_data <= 16'h0000;
            12'd2173 : o_data <= 16'h0000;
            12'd2174 : o_data <= 16'h0000;
            12'd2175 : o_data <= 16'h0000;
            12'd2176 : o_data <= 16'h0000;
            12'd2177 : o_data <= 16'h0000;
            12'd2178 : o_data <= 16'h0000;
            12'd2179 : o_data <= 16'h0000;
            12'd2180 : o_data <= 16'h0000;
            12'd2181 : o_data <= 16'h0000;
            12'd2182 : o_data <= 16'h0000;
            12'd2183 : o_data <= 16'h0000;
            12'd2184 : o_data <= 16'h0000;
            12'd2185 : o_data <= 16'h0000;
            12'd2186 : o_data <= 16'h0000;
            12'd2187 : o_data <= 16'h0000;
            12'd2188 : o_data <= 16'h0000;
            12'd2189 : o_data <= 16'h0000;
            12'd2190 : o_data <= 16'h0000;
            12'd2191 : o_data <= 16'h0000;
            12'd2192 : o_data <= 16'h0000;
            12'd2193 : o_data <= 16'h0000;
            12'd2194 : o_data <= 16'h0000;
            12'd2195 : o_data <= 16'h0000;
            12'd2196 : o_data <= 16'h0000;
            12'd2197 : o_data <= 16'h0000;
            12'd2198 : o_data <= 16'h0000;
            12'd2199 : o_data <= 16'h0000;
            12'd2200 : o_data <= 16'h0000;
            12'd2201 : o_data <= 16'h0000;
            12'd2202 : o_data <= 16'h0000;
            12'd2203 : o_data <= 16'h0000;
            12'd2204 : o_data <= 16'h0000;
            12'd2205 : o_data <= 16'h0000;
            12'd2206 : o_data <= 16'h0000;
            12'd2207 : o_data <= 16'h0000;
            12'd2208 : o_data <= 16'h0000;
            12'd2209 : o_data <= 16'h0000;
            12'd2210 : o_data <= 16'h0000;
            12'd2211 : o_data <= 16'h0000;
            12'd2212 : o_data <= 16'h0000;
            12'd2213 : o_data <= 16'h0000;
            12'd2214 : o_data <= 16'h0000;
            12'd2215 : o_data <= 16'h0000;
            12'd2216 : o_data <= 16'h0000;
            12'd2217 : o_data <= 16'h0000;
            12'd2218 : o_data <= 16'h0000;
            12'd2219 : o_data <= 16'h0000;
            12'd2220 : o_data <= 16'h0000;
            12'd2221 : o_data <= 16'h0000;
            12'd2222 : o_data <= 16'h0000;
            12'd2223 : o_data <= 16'h0000;
            12'd2224 : o_data <= 16'h0000;
            12'd2225 : o_data <= 16'h0000;
            12'd2226 : o_data <= 16'h0000;
            12'd2227 : o_data <= 16'h0000;
            12'd2228 : o_data <= 16'h0000;
            12'd2229 : o_data <= 16'h0000;
            12'd2230 : o_data <= 16'h0000;
            12'd2231 : o_data <= 16'h0000;
            12'd2232 : o_data <= 16'h0000;
            12'd2233 : o_data <= 16'h0000;
            12'd2234 : o_data <= 16'h0000;
            12'd2235 : o_data <= 16'h0000;
            12'd2236 : o_data <= 16'h0000;
            12'd2237 : o_data <= 16'h0000;
            12'd2238 : o_data <= 16'h0000;
            12'd2239 : o_data <= 16'h0000;
            12'd2240 : o_data <= 16'h0000;
            12'd2241 : o_data <= 16'h0000;
            12'd2242 : o_data <= 16'h0000;
            12'd2243 : o_data <= 16'h0000;
            12'd2244 : o_data <= 16'h0000;
            12'd2245 : o_data <= 16'h0000;
            12'd2246 : o_data <= 16'h0000;
            12'd2247 : o_data <= 16'h0000;
            12'd2248 : o_data <= 16'h0000;
            12'd2249 : o_data <= 16'h0000;
            12'd2250 : o_data <= 16'h0000;
            12'd2251 : o_data <= 16'h0000;
            12'd2252 : o_data <= 16'h0000;
            12'd2253 : o_data <= 16'h0000;
            12'd2254 : o_data <= 16'h0000;
            12'd2255 : o_data <= 16'h0000;
            12'd2256 : o_data <= 16'h0000;
            12'd2257 : o_data <= 16'h0000;
            12'd2258 : o_data <= 16'h0000;
            12'd2259 : o_data <= 16'h0000;
            12'd2260 : o_data <= 16'h0000;
            12'd2261 : o_data <= 16'h0000;
            12'd2262 : o_data <= 16'h0000;
            12'd2263 : o_data <= 16'h0000;
            12'd2264 : o_data <= 16'h0000;
            12'd2265 : o_data <= 16'h0000;
            12'd2266 : o_data <= 16'h0000;
            12'd2267 : o_data <= 16'h0000;
            12'd2268 : o_data <= 16'h0000;
            12'd2269 : o_data <= 16'h0000;
            12'd2270 : o_data <= 16'h0000;
            12'd2271 : o_data <= 16'h0000;
            12'd2272 : o_data <= 16'h0000;
            12'd2273 : o_data <= 16'h0000;
            12'd2274 : o_data <= 16'h0000;
            12'd2275 : o_data <= 16'h0000;
            12'd2276 : o_data <= 16'h0000;
            12'd2277 : o_data <= 16'h0000;
            12'd2278 : o_data <= 16'h0000;
            12'd2279 : o_data <= 16'h0000;
            12'd2280 : o_data <= 16'h0000;
            12'd2281 : o_data <= 16'h0000;
            12'd2282 : o_data <= 16'h0000;
            12'd2283 : o_data <= 16'h0000;
            12'd2284 : o_data <= 16'h0000;
            12'd2285 : o_data <= 16'h0000;
            12'd2286 : o_data <= 16'h0000;
            12'd2287 : o_data <= 16'h0000;
            12'd2288 : o_data <= 16'h0000;
            12'd2289 : o_data <= 16'h0000;
            12'd2290 : o_data <= 16'h0000;
            12'd2291 : o_data <= 16'h0000;
            12'd2292 : o_data <= 16'h0000;
            12'd2293 : o_data <= 16'h0000;
            12'd2294 : o_data <= 16'h0000;
            12'd2295 : o_data <= 16'h0000;
            12'd2296 : o_data <= 16'h0000;
            12'd2297 : o_data <= 16'h0000;
            12'd2298 : o_data <= 16'h0000;
            12'd2299 : o_data <= 16'h0000;
            12'd2300 : o_data <= 16'h0000;
            12'd2301 : o_data <= 16'h0000;
            12'd2302 : o_data <= 16'h0000;
            12'd2303 : o_data <= 16'h0000;
            default : o_data <= 16'd0;
        endcase
    end

endmodule
